magic
tech sky130A
magscale 1 2
timestamp 1624067825
<< obsli1 >>
rect 1104 1513 78844 77809
<< obsm1 >>
rect 106 1368 79842 78600
<< metal2 >>
rect 110 79200 166 80800
rect 386 79200 442 80800
rect 754 79200 810 80800
rect 1030 79200 1086 80800
rect 1398 79200 1454 80800
rect 1674 79200 1730 80800
rect 2042 79200 2098 80800
rect 2410 79200 2466 80800
rect 2686 79200 2742 80800
rect 3054 79200 3110 80800
rect 3330 79200 3386 80800
rect 3698 79200 3754 80800
rect 3974 79200 4030 80800
rect 4342 79200 4398 80800
rect 4710 79200 4766 80800
rect 4986 79200 5042 80800
rect 5354 79200 5410 80800
rect 5630 79200 5686 80800
rect 5998 79200 6054 80800
rect 6366 79200 6422 80800
rect 6642 79200 6698 80800
rect 7010 79200 7066 80800
rect 7286 79200 7342 80800
rect 7654 79200 7710 80800
rect 7930 79200 7986 80800
rect 8298 79200 8354 80800
rect 8666 79200 8722 80800
rect 8942 79200 8998 80800
rect 9310 79200 9366 80800
rect 9586 79200 9642 80800
rect 9954 79200 10010 80800
rect 10230 79200 10286 80800
rect 10598 79200 10654 80800
rect 10966 79200 11022 80800
rect 11242 79200 11298 80800
rect 11610 79200 11666 80800
rect 11886 79200 11942 80800
rect 12254 79200 12310 80800
rect 12622 79200 12678 80800
rect 12898 79200 12954 80800
rect 13266 79200 13322 80800
rect 13542 79200 13598 80800
rect 13910 79200 13966 80800
rect 14186 79200 14242 80800
rect 14554 79200 14610 80800
rect 14922 79200 14978 80800
rect 15198 79200 15254 80800
rect 15566 79200 15622 80800
rect 15842 79200 15898 80800
rect 16210 79200 16266 80800
rect 16578 79200 16634 80800
rect 16854 79200 16910 80800
rect 17222 79200 17278 80800
rect 17498 79200 17554 80800
rect 17866 79200 17922 80800
rect 18142 79200 18198 80800
rect 18510 79200 18566 80800
rect 18878 79200 18934 80800
rect 19154 79200 19210 80800
rect 19522 79200 19578 80800
rect 19798 79200 19854 80800
rect 20166 79200 20222 80800
rect 20442 79200 20498 80800
rect 20810 79200 20866 80800
rect 21178 79200 21234 80800
rect 21454 79200 21510 80800
rect 21822 79200 21878 80800
rect 22098 79200 22154 80800
rect 22466 79200 22522 80800
rect 22834 79200 22890 80800
rect 23110 79200 23166 80800
rect 23478 79200 23534 80800
rect 23754 79200 23810 80800
rect 24122 79200 24178 80800
rect 24398 79200 24454 80800
rect 24766 79200 24822 80800
rect 25134 79200 25190 80800
rect 25410 79200 25466 80800
rect 25778 79200 25834 80800
rect 26054 79200 26110 80800
rect 26422 79200 26478 80800
rect 26790 79200 26846 80800
rect 27066 79200 27122 80800
rect 27434 79200 27490 80800
rect 27710 79200 27766 80800
rect 28078 79200 28134 80800
rect 28354 79200 28410 80800
rect 28722 79200 28778 80800
rect 29090 79200 29146 80800
rect 29366 79200 29422 80800
rect 29734 79200 29790 80800
rect 30010 79200 30066 80800
rect 30378 79200 30434 80800
rect 30654 79200 30710 80800
rect 31022 79200 31078 80800
rect 31390 79200 31446 80800
rect 31666 79200 31722 80800
rect 32034 79200 32090 80800
rect 32310 79200 32366 80800
rect 32678 79200 32734 80800
rect 33046 79200 33102 80800
rect 33322 79200 33378 80800
rect 33690 79200 33746 80800
rect 33966 79200 34022 80800
rect 34334 79200 34390 80800
rect 34610 79200 34666 80800
rect 34978 79200 35034 80800
rect 35346 79200 35402 80800
rect 35622 79200 35678 80800
rect 35990 79200 36046 80800
rect 36266 79200 36322 80800
rect 36634 79200 36690 80800
rect 36910 79200 36966 80800
rect 37278 79200 37334 80800
rect 37646 79200 37702 80800
rect 37922 79200 37978 80800
rect 38290 79200 38346 80800
rect 38566 79200 38622 80800
rect 38934 79200 38990 80800
rect 39302 79200 39358 80800
rect 39578 79200 39634 80800
rect 39946 79200 40002 80800
rect 40222 79200 40278 80800
rect 40590 79200 40646 80800
rect 40866 79200 40922 80800
rect 41234 79200 41290 80800
rect 41602 79200 41658 80800
rect 41878 79200 41934 80800
rect 42246 79200 42302 80800
rect 42522 79200 42578 80800
rect 42890 79200 42946 80800
rect 43258 79200 43314 80800
rect 43534 79200 43590 80800
rect 43902 79200 43958 80800
rect 44178 79200 44234 80800
rect 44546 79200 44602 80800
rect 44822 79200 44878 80800
rect 45190 79200 45246 80800
rect 45558 79200 45614 80800
rect 45834 79200 45890 80800
rect 46202 79200 46258 80800
rect 46478 79200 46534 80800
rect 46846 79200 46902 80800
rect 47122 79200 47178 80800
rect 47490 79200 47546 80800
rect 47858 79200 47914 80800
rect 48134 79200 48190 80800
rect 48502 79200 48558 80800
rect 48778 79200 48834 80800
rect 49146 79200 49202 80800
rect 49514 79200 49570 80800
rect 49790 79200 49846 80800
rect 50158 79200 50214 80800
rect 50434 79200 50490 80800
rect 50802 79200 50858 80800
rect 51078 79200 51134 80800
rect 51446 79200 51502 80800
rect 51814 79200 51870 80800
rect 52090 79200 52146 80800
rect 52458 79200 52514 80800
rect 52734 79200 52790 80800
rect 53102 79200 53158 80800
rect 53470 79200 53526 80800
rect 53746 79200 53802 80800
rect 54114 79200 54170 80800
rect 54390 79200 54446 80800
rect 54758 79200 54814 80800
rect 55034 79200 55090 80800
rect 55402 79200 55458 80800
rect 55770 79200 55826 80800
rect 56046 79200 56102 80800
rect 56414 79200 56470 80800
rect 56690 79200 56746 80800
rect 57058 79200 57114 80800
rect 57334 79200 57390 80800
rect 57702 79200 57758 80800
rect 58070 79200 58126 80800
rect 58346 79200 58402 80800
rect 58714 79200 58770 80800
rect 58990 79200 59046 80800
rect 59358 79200 59414 80800
rect 59726 79200 59782 80800
rect 60002 79200 60058 80800
rect 60370 79200 60426 80800
rect 60646 79200 60702 80800
rect 61014 79200 61070 80800
rect 61290 79200 61346 80800
rect 61658 79200 61714 80800
rect 62026 79200 62082 80800
rect 62302 79200 62358 80800
rect 62670 79200 62726 80800
rect 62946 79200 63002 80800
rect 63314 79200 63370 80800
rect 63590 79200 63646 80800
rect 63958 79200 64014 80800
rect 64326 79200 64382 80800
rect 64602 79200 64658 80800
rect 64970 79200 65026 80800
rect 65246 79200 65302 80800
rect 65614 79200 65670 80800
rect 65982 79200 66038 80800
rect 66258 79200 66314 80800
rect 66626 79200 66682 80800
rect 66902 79200 66958 80800
rect 67270 79200 67326 80800
rect 67546 79200 67602 80800
rect 67914 79200 67970 80800
rect 68282 79200 68338 80800
rect 68558 79200 68614 80800
rect 68926 79200 68982 80800
rect 69202 79200 69258 80800
rect 69570 79200 69626 80800
rect 69938 79200 69994 80800
rect 70214 79200 70270 80800
rect 70582 79200 70638 80800
rect 70858 79200 70914 80800
rect 71226 79200 71282 80800
rect 71502 79200 71558 80800
rect 71870 79200 71926 80800
rect 72238 79200 72294 80800
rect 72514 79200 72570 80800
rect 72882 79200 72938 80800
rect 73158 79200 73214 80800
rect 73526 79200 73582 80800
rect 73802 79200 73858 80800
rect 74170 79200 74226 80800
rect 74538 79200 74594 80800
rect 74814 79200 74870 80800
rect 75182 79200 75238 80800
rect 75458 79200 75514 80800
rect 75826 79200 75882 80800
rect 76194 79200 76250 80800
rect 76470 79200 76526 80800
rect 76838 79200 76894 80800
rect 77114 79200 77170 80800
rect 77482 79200 77538 80800
rect 77758 79200 77814 80800
rect 78126 79200 78182 80800
rect 78494 79200 78550 80800
rect 78770 79200 78826 80800
rect 79138 79200 79194 80800
rect 79414 79200 79470 80800
rect 79782 79200 79838 80800
rect 294 -800 350 800
rect 846 -800 902 800
rect 1490 -800 1546 800
rect 2134 -800 2190 800
rect 2778 -800 2834 800
rect 3330 -800 3386 800
rect 3974 -800 4030 800
rect 4618 -800 4674 800
rect 5262 -800 5318 800
rect 5906 -800 5962 800
rect 6458 -800 6514 800
rect 7102 -800 7158 800
rect 7746 -800 7802 800
rect 8390 -800 8446 800
rect 9034 -800 9090 800
rect 9586 -800 9642 800
rect 10230 -800 10286 800
rect 10874 -800 10930 800
rect 11518 -800 11574 800
rect 12162 -800 12218 800
rect 12714 -800 12770 800
rect 13358 -800 13414 800
rect 14002 -800 14058 800
rect 14646 -800 14702 800
rect 15290 -800 15346 800
rect 15842 -800 15898 800
rect 16486 -800 16542 800
rect 17130 -800 17186 800
rect 17774 -800 17830 800
rect 18418 -800 18474 800
rect 18970 -800 19026 800
rect 19614 -800 19670 800
rect 20258 -800 20314 800
rect 20902 -800 20958 800
rect 21546 -800 21602 800
rect 22098 -800 22154 800
rect 22742 -800 22798 800
rect 23386 -800 23442 800
rect 24030 -800 24086 800
rect 24674 -800 24730 800
rect 25226 -800 25282 800
rect 25870 -800 25926 800
rect 26514 -800 26570 800
rect 27158 -800 27214 800
rect 27802 -800 27858 800
rect 28354 -800 28410 800
rect 28998 -800 29054 800
rect 29642 -800 29698 800
rect 30286 -800 30342 800
rect 30930 -800 30986 800
rect 31482 -800 31538 800
rect 32126 -800 32182 800
rect 32770 -800 32826 800
rect 33414 -800 33470 800
rect 34058 -800 34114 800
rect 34610 -800 34666 800
rect 35254 -800 35310 800
rect 35898 -800 35954 800
rect 36542 -800 36598 800
rect 37186 -800 37242 800
rect 37738 -800 37794 800
rect 38382 -800 38438 800
rect 39026 -800 39082 800
rect 39670 -800 39726 800
rect 40314 -800 40370 800
rect 40866 -800 40922 800
rect 41510 -800 41566 800
rect 42154 -800 42210 800
rect 42798 -800 42854 800
rect 43350 -800 43406 800
rect 43994 -800 44050 800
rect 44638 -800 44694 800
rect 45282 -800 45338 800
rect 45926 -800 45982 800
rect 46478 -800 46534 800
rect 47122 -800 47178 800
rect 47766 -800 47822 800
rect 48410 -800 48466 800
rect 49054 -800 49110 800
rect 49606 -800 49662 800
rect 50250 -800 50306 800
rect 50894 -800 50950 800
rect 51538 -800 51594 800
rect 52182 -800 52238 800
rect 52734 -800 52790 800
rect 53378 -800 53434 800
rect 54022 -800 54078 800
rect 54666 -800 54722 800
rect 55310 -800 55366 800
rect 55862 -800 55918 800
rect 56506 -800 56562 800
rect 57150 -800 57206 800
rect 57794 -800 57850 800
rect 58438 -800 58494 800
rect 58990 -800 59046 800
rect 59634 -800 59690 800
rect 60278 -800 60334 800
rect 60922 -800 60978 800
rect 61566 -800 61622 800
rect 62118 -800 62174 800
rect 62762 -800 62818 800
rect 63406 -800 63462 800
rect 64050 -800 64106 800
rect 64694 -800 64750 800
rect 65246 -800 65302 800
rect 65890 -800 65946 800
rect 66534 -800 66590 800
rect 67178 -800 67234 800
rect 67822 -800 67878 800
rect 68374 -800 68430 800
rect 69018 -800 69074 800
rect 69662 -800 69718 800
rect 70306 -800 70362 800
rect 70950 -800 71006 800
rect 71502 -800 71558 800
rect 72146 -800 72202 800
rect 72790 -800 72846 800
rect 73434 -800 73490 800
rect 74078 -800 74134 800
rect 74630 -800 74686 800
rect 75274 -800 75330 800
rect 75918 -800 75974 800
rect 76562 -800 76618 800
rect 77206 -800 77262 800
rect 77758 -800 77814 800
rect 78402 -800 78458 800
rect 79046 -800 79102 800
rect 79690 -800 79746 800
<< obsm2 >>
rect 222 79144 330 79801
rect 498 79144 698 79801
rect 866 79144 974 79801
rect 1142 79144 1342 79801
rect 1510 79144 1618 79801
rect 1786 79144 1986 79801
rect 2154 79144 2354 79801
rect 2522 79144 2630 79801
rect 2798 79144 2998 79801
rect 3166 79144 3274 79801
rect 3442 79144 3642 79801
rect 3810 79144 3918 79801
rect 4086 79144 4286 79801
rect 4454 79144 4654 79801
rect 4822 79144 4930 79801
rect 5098 79144 5298 79801
rect 5466 79144 5574 79801
rect 5742 79144 5942 79801
rect 6110 79144 6310 79801
rect 6478 79144 6586 79801
rect 6754 79144 6954 79801
rect 7122 79144 7230 79801
rect 7398 79144 7598 79801
rect 7766 79144 7874 79801
rect 8042 79144 8242 79801
rect 8410 79144 8610 79801
rect 8778 79144 8886 79801
rect 9054 79144 9254 79801
rect 9422 79144 9530 79801
rect 9698 79144 9898 79801
rect 10066 79144 10174 79801
rect 10342 79144 10542 79801
rect 10710 79144 10910 79801
rect 11078 79144 11186 79801
rect 11354 79144 11554 79801
rect 11722 79144 11830 79801
rect 11998 79144 12198 79801
rect 12366 79144 12566 79801
rect 12734 79144 12842 79801
rect 13010 79144 13210 79801
rect 13378 79144 13486 79801
rect 13654 79144 13854 79801
rect 14022 79144 14130 79801
rect 14298 79144 14498 79801
rect 14666 79144 14866 79801
rect 15034 79144 15142 79801
rect 15310 79144 15510 79801
rect 15678 79144 15786 79801
rect 15954 79144 16154 79801
rect 16322 79144 16522 79801
rect 16690 79144 16798 79801
rect 16966 79144 17166 79801
rect 17334 79144 17442 79801
rect 17610 79144 17810 79801
rect 17978 79144 18086 79801
rect 18254 79144 18454 79801
rect 18622 79144 18822 79801
rect 18990 79144 19098 79801
rect 19266 79144 19466 79801
rect 19634 79144 19742 79801
rect 19910 79144 20110 79801
rect 20278 79144 20386 79801
rect 20554 79144 20754 79801
rect 20922 79144 21122 79801
rect 21290 79144 21398 79801
rect 21566 79144 21766 79801
rect 21934 79144 22042 79801
rect 22210 79144 22410 79801
rect 22578 79144 22778 79801
rect 22946 79144 23054 79801
rect 23222 79144 23422 79801
rect 23590 79144 23698 79801
rect 23866 79144 24066 79801
rect 24234 79144 24342 79801
rect 24510 79144 24710 79801
rect 24878 79144 25078 79801
rect 25246 79144 25354 79801
rect 25522 79144 25722 79801
rect 25890 79144 25998 79801
rect 26166 79144 26366 79801
rect 26534 79144 26734 79801
rect 26902 79144 27010 79801
rect 27178 79144 27378 79801
rect 27546 79144 27654 79801
rect 27822 79144 28022 79801
rect 28190 79144 28298 79801
rect 28466 79144 28666 79801
rect 28834 79144 29034 79801
rect 29202 79144 29310 79801
rect 29478 79144 29678 79801
rect 29846 79144 29954 79801
rect 30122 79144 30322 79801
rect 30490 79144 30598 79801
rect 30766 79144 30966 79801
rect 31134 79144 31334 79801
rect 31502 79144 31610 79801
rect 31778 79144 31978 79801
rect 32146 79144 32254 79801
rect 32422 79144 32622 79801
rect 32790 79144 32990 79801
rect 33158 79144 33266 79801
rect 33434 79144 33634 79801
rect 33802 79144 33910 79801
rect 34078 79144 34278 79801
rect 34446 79144 34554 79801
rect 34722 79144 34922 79801
rect 35090 79144 35290 79801
rect 35458 79144 35566 79801
rect 35734 79144 35934 79801
rect 36102 79144 36210 79801
rect 36378 79144 36578 79801
rect 36746 79144 36854 79801
rect 37022 79144 37222 79801
rect 37390 79144 37590 79801
rect 37758 79144 37866 79801
rect 38034 79144 38234 79801
rect 38402 79144 38510 79801
rect 38678 79144 38878 79801
rect 39046 79144 39246 79801
rect 39414 79144 39522 79801
rect 39690 79144 39890 79801
rect 40058 79144 40166 79801
rect 40334 79144 40534 79801
rect 40702 79144 40810 79801
rect 40978 79144 41178 79801
rect 41346 79144 41546 79801
rect 41714 79144 41822 79801
rect 41990 79144 42190 79801
rect 42358 79144 42466 79801
rect 42634 79144 42834 79801
rect 43002 79144 43202 79801
rect 43370 79144 43478 79801
rect 43646 79144 43846 79801
rect 44014 79144 44122 79801
rect 44290 79144 44490 79801
rect 44658 79144 44766 79801
rect 44934 79144 45134 79801
rect 45302 79144 45502 79801
rect 45670 79144 45778 79801
rect 45946 79144 46146 79801
rect 46314 79144 46422 79801
rect 46590 79144 46790 79801
rect 46958 79144 47066 79801
rect 47234 79144 47434 79801
rect 47602 79144 47802 79801
rect 47970 79144 48078 79801
rect 48246 79144 48446 79801
rect 48614 79144 48722 79801
rect 48890 79144 49090 79801
rect 49258 79144 49458 79801
rect 49626 79144 49734 79801
rect 49902 79144 50102 79801
rect 50270 79144 50378 79801
rect 50546 79144 50746 79801
rect 50914 79144 51022 79801
rect 51190 79144 51390 79801
rect 51558 79144 51758 79801
rect 51926 79144 52034 79801
rect 52202 79144 52402 79801
rect 52570 79144 52678 79801
rect 52846 79144 53046 79801
rect 53214 79144 53414 79801
rect 53582 79144 53690 79801
rect 53858 79144 54058 79801
rect 54226 79144 54334 79801
rect 54502 79144 54702 79801
rect 54870 79144 54978 79801
rect 55146 79144 55346 79801
rect 55514 79144 55714 79801
rect 55882 79144 55990 79801
rect 56158 79144 56358 79801
rect 56526 79144 56634 79801
rect 56802 79144 57002 79801
rect 57170 79144 57278 79801
rect 57446 79144 57646 79801
rect 57814 79144 58014 79801
rect 58182 79144 58290 79801
rect 58458 79144 58658 79801
rect 58826 79144 58934 79801
rect 59102 79144 59302 79801
rect 59470 79144 59670 79801
rect 59838 79144 59946 79801
rect 60114 79144 60314 79801
rect 60482 79144 60590 79801
rect 60758 79144 60958 79801
rect 61126 79144 61234 79801
rect 61402 79144 61602 79801
rect 61770 79144 61970 79801
rect 62138 79144 62246 79801
rect 62414 79144 62614 79801
rect 62782 79144 62890 79801
rect 63058 79144 63258 79801
rect 63426 79144 63534 79801
rect 63702 79144 63902 79801
rect 64070 79144 64270 79801
rect 64438 79144 64546 79801
rect 64714 79144 64914 79801
rect 65082 79144 65190 79801
rect 65358 79144 65558 79801
rect 65726 79144 65926 79801
rect 66094 79144 66202 79801
rect 66370 79144 66570 79801
rect 66738 79144 66846 79801
rect 67014 79144 67214 79801
rect 67382 79144 67490 79801
rect 67658 79144 67858 79801
rect 68026 79144 68226 79801
rect 68394 79144 68502 79801
rect 68670 79144 68870 79801
rect 69038 79144 69146 79801
rect 69314 79144 69514 79801
rect 69682 79144 69882 79801
rect 70050 79144 70158 79801
rect 70326 79144 70526 79801
rect 70694 79144 70802 79801
rect 70970 79144 71170 79801
rect 71338 79144 71446 79801
rect 71614 79144 71814 79801
rect 71982 79144 72182 79801
rect 72350 79144 72458 79801
rect 72626 79144 72826 79801
rect 72994 79144 73102 79801
rect 73270 79144 73470 79801
rect 73638 79144 73746 79801
rect 73914 79144 74114 79801
rect 74282 79144 74482 79801
rect 74650 79144 74758 79801
rect 74926 79144 75126 79801
rect 75294 79144 75402 79801
rect 75570 79144 75770 79801
rect 75938 79144 76138 79801
rect 76306 79144 76414 79801
rect 76582 79144 76782 79801
rect 76950 79144 77058 79801
rect 77226 79144 77426 79801
rect 77594 79144 77702 79801
rect 77870 79144 78070 79801
rect 78238 79144 78438 79801
rect 78606 79144 78714 79801
rect 78882 79144 79082 79801
rect 79250 79144 79358 79801
rect 79526 79144 79726 79801
rect 112 856 79836 79144
rect 112 303 238 856
rect 406 303 790 856
rect 958 303 1434 856
rect 1602 303 2078 856
rect 2246 303 2722 856
rect 2890 303 3274 856
rect 3442 303 3918 856
rect 4086 303 4562 856
rect 4730 303 5206 856
rect 5374 303 5850 856
rect 6018 303 6402 856
rect 6570 303 7046 856
rect 7214 303 7690 856
rect 7858 303 8334 856
rect 8502 303 8978 856
rect 9146 303 9530 856
rect 9698 303 10174 856
rect 10342 303 10818 856
rect 10986 303 11462 856
rect 11630 303 12106 856
rect 12274 303 12658 856
rect 12826 303 13302 856
rect 13470 303 13946 856
rect 14114 303 14590 856
rect 14758 303 15234 856
rect 15402 303 15786 856
rect 15954 303 16430 856
rect 16598 303 17074 856
rect 17242 303 17718 856
rect 17886 303 18362 856
rect 18530 303 18914 856
rect 19082 303 19558 856
rect 19726 303 20202 856
rect 20370 303 20846 856
rect 21014 303 21490 856
rect 21658 303 22042 856
rect 22210 303 22686 856
rect 22854 303 23330 856
rect 23498 303 23974 856
rect 24142 303 24618 856
rect 24786 303 25170 856
rect 25338 303 25814 856
rect 25982 303 26458 856
rect 26626 303 27102 856
rect 27270 303 27746 856
rect 27914 303 28298 856
rect 28466 303 28942 856
rect 29110 303 29586 856
rect 29754 303 30230 856
rect 30398 303 30874 856
rect 31042 303 31426 856
rect 31594 303 32070 856
rect 32238 303 32714 856
rect 32882 303 33358 856
rect 33526 303 34002 856
rect 34170 303 34554 856
rect 34722 303 35198 856
rect 35366 303 35842 856
rect 36010 303 36486 856
rect 36654 303 37130 856
rect 37298 303 37682 856
rect 37850 303 38326 856
rect 38494 303 38970 856
rect 39138 303 39614 856
rect 39782 303 40258 856
rect 40426 303 40810 856
rect 40978 303 41454 856
rect 41622 303 42098 856
rect 42266 303 42742 856
rect 42910 303 43294 856
rect 43462 303 43938 856
rect 44106 303 44582 856
rect 44750 303 45226 856
rect 45394 303 45870 856
rect 46038 303 46422 856
rect 46590 303 47066 856
rect 47234 303 47710 856
rect 47878 303 48354 856
rect 48522 303 48998 856
rect 49166 303 49550 856
rect 49718 303 50194 856
rect 50362 303 50838 856
rect 51006 303 51482 856
rect 51650 303 52126 856
rect 52294 303 52678 856
rect 52846 303 53322 856
rect 53490 303 53966 856
rect 54134 303 54610 856
rect 54778 303 55254 856
rect 55422 303 55806 856
rect 55974 303 56450 856
rect 56618 303 57094 856
rect 57262 303 57738 856
rect 57906 303 58382 856
rect 58550 303 58934 856
rect 59102 303 59578 856
rect 59746 303 60222 856
rect 60390 303 60866 856
rect 61034 303 61510 856
rect 61678 303 62062 856
rect 62230 303 62706 856
rect 62874 303 63350 856
rect 63518 303 63994 856
rect 64162 303 64638 856
rect 64806 303 65190 856
rect 65358 303 65834 856
rect 66002 303 66478 856
rect 66646 303 67122 856
rect 67290 303 67766 856
rect 67934 303 68318 856
rect 68486 303 68962 856
rect 69130 303 69606 856
rect 69774 303 70250 856
rect 70418 303 70894 856
rect 71062 303 71446 856
rect 71614 303 72090 856
rect 72258 303 72734 856
rect 72902 303 73378 856
rect 73546 303 74022 856
rect 74190 303 74574 856
rect 74742 303 75218 856
rect 75386 303 75862 856
rect 76030 303 76506 856
rect 76674 303 77150 856
rect 77318 303 77702 856
rect 77870 303 78346 856
rect 78514 303 78990 856
rect 79158 303 79634 856
rect 79802 303 79836 856
<< metal3 >>
rect -800 79704 800 79824
rect 79200 79568 80800 79688
rect -800 79296 800 79416
rect -800 78888 800 79008
rect 79200 78888 80800 79008
rect -800 78480 800 78600
rect 79200 78344 80800 78464
rect -800 78072 800 78192
rect -800 77664 800 77784
rect 79200 77664 80800 77784
rect -800 77256 800 77376
rect 79200 77120 80800 77240
rect -800 76848 800 76968
rect -800 76440 800 76560
rect 79200 76440 80800 76560
rect -800 76032 800 76152
rect -800 75624 800 75744
rect 79200 75760 80800 75880
rect -800 75216 800 75336
rect 79200 75216 80800 75336
rect -800 74808 800 74928
rect -800 74400 800 74520
rect 79200 74536 80800 74656
rect -800 73992 800 74112
rect 79200 73992 80800 74112
rect -800 73584 800 73704
rect -800 73176 800 73296
rect 79200 73312 80800 73432
rect -800 72768 800 72888
rect 79200 72632 80800 72752
rect -800 72360 800 72480
rect -800 71952 800 72072
rect 79200 72088 80800 72208
rect -800 71544 800 71664
rect 79200 71408 80800 71528
rect -800 71136 800 71256
rect -800 70864 800 70984
rect 79200 70864 80800 70984
rect -800 70456 800 70576
rect -800 70048 800 70168
rect 79200 70184 80800 70304
rect -800 69640 800 69760
rect 79200 69504 80800 69624
rect -800 69232 800 69352
rect -800 68824 800 68944
rect 79200 68960 80800 69080
rect -800 68416 800 68536
rect 79200 68280 80800 68400
rect -800 68008 800 68128
rect -800 67600 800 67720
rect 79200 67736 80800 67856
rect -800 67192 800 67312
rect 79200 67056 80800 67176
rect -800 66784 800 66904
rect -800 66376 800 66496
rect 79200 66376 80800 66496
rect -800 65968 800 66088
rect 79200 65832 80800 65952
rect -800 65560 800 65680
rect -800 65152 800 65272
rect 79200 65152 80800 65272
rect -800 64744 800 64864
rect 79200 64608 80800 64728
rect -800 64336 800 64456
rect -800 63928 800 64048
rect 79200 63928 80800 64048
rect -800 63520 800 63640
rect -800 63112 800 63232
rect 79200 63248 80800 63368
rect -800 62704 800 62824
rect 79200 62704 80800 62824
rect -800 62296 800 62416
rect -800 62024 800 62144
rect 79200 62024 80800 62144
rect -800 61616 800 61736
rect 79200 61480 80800 61600
rect -800 61208 800 61328
rect -800 60800 800 60920
rect 79200 60800 80800 60920
rect -800 60392 800 60512
rect 79200 60256 80800 60376
rect -800 59984 800 60104
rect -800 59576 800 59696
rect 79200 59576 80800 59696
rect -800 59168 800 59288
rect -800 58760 800 58880
rect 79200 58896 80800 59016
rect -800 58352 800 58472
rect 79200 58352 80800 58472
rect -800 57944 800 58064
rect -800 57536 800 57656
rect 79200 57672 80800 57792
rect -800 57128 800 57248
rect 79200 57128 80800 57248
rect -800 56720 800 56840
rect -800 56312 800 56432
rect 79200 56448 80800 56568
rect -800 55904 800 56024
rect 79200 55768 80800 55888
rect -800 55496 800 55616
rect -800 55088 800 55208
rect 79200 55224 80800 55344
rect -800 54680 800 54800
rect 79200 54544 80800 54664
rect -800 54272 800 54392
rect -800 53864 800 53984
rect 79200 54000 80800 54120
rect -800 53456 800 53576
rect -800 53184 800 53304
rect 79200 53320 80800 53440
rect -800 52776 800 52896
rect 79200 52640 80800 52760
rect -800 52368 800 52488
rect -800 51960 800 52080
rect 79200 52096 80800 52216
rect -800 51552 800 51672
rect 79200 51416 80800 51536
rect -800 51144 800 51264
rect -800 50736 800 50856
rect 79200 50872 80800 50992
rect -800 50328 800 50448
rect 79200 50192 80800 50312
rect -800 49920 800 50040
rect -800 49512 800 49632
rect 79200 49512 80800 49632
rect -800 49104 800 49224
rect 79200 48968 80800 49088
rect -800 48696 800 48816
rect -800 48288 800 48408
rect 79200 48288 80800 48408
rect -800 47880 800 48000
rect 79200 47744 80800 47864
rect -800 47472 800 47592
rect -800 47064 800 47184
rect 79200 47064 80800 47184
rect -800 46656 800 46776
rect -800 46248 800 46368
rect 79200 46384 80800 46504
rect -800 45840 800 45960
rect 79200 45840 80800 45960
rect -800 45432 800 45552
rect -800 45024 800 45144
rect 79200 45160 80800 45280
rect -800 44616 800 44736
rect 79200 44616 80800 44736
rect -800 44344 800 44464
rect -800 43936 800 44056
rect 79200 43936 80800 44056
rect -800 43528 800 43648
rect -800 43120 800 43240
rect 79200 43256 80800 43376
rect -800 42712 800 42832
rect 79200 42712 80800 42832
rect -800 42304 800 42424
rect -800 41896 800 42016
rect 79200 42032 80800 42152
rect -800 41488 800 41608
rect 79200 41488 80800 41608
rect -800 41080 800 41200
rect -800 40672 800 40792
rect 79200 40808 80800 40928
rect -800 40264 800 40384
rect 79200 40264 80800 40384
rect -800 39856 800 39976
rect -800 39448 800 39568
rect 79200 39584 80800 39704
rect -800 39040 800 39160
rect 79200 38904 80800 39024
rect -800 38632 800 38752
rect -800 38224 800 38344
rect 79200 38360 80800 38480
rect -800 37816 800 37936
rect 79200 37680 80800 37800
rect -800 37408 800 37528
rect -800 37000 800 37120
rect 79200 37136 80800 37256
rect -800 36592 800 36712
rect 79200 36456 80800 36576
rect -800 36184 800 36304
rect -800 35776 800 35896
rect 79200 35776 80800 35896
rect -800 35504 800 35624
rect -800 35096 800 35216
rect 79200 35232 80800 35352
rect -800 34688 800 34808
rect 79200 34552 80800 34672
rect -800 34280 800 34400
rect -800 33872 800 33992
rect 79200 34008 80800 34128
rect -800 33464 800 33584
rect 79200 33328 80800 33448
rect -800 33056 800 33176
rect -800 32648 800 32768
rect 79200 32648 80800 32768
rect -800 32240 800 32360
rect 79200 32104 80800 32224
rect -800 31832 800 31952
rect -800 31424 800 31544
rect 79200 31424 80800 31544
rect -800 31016 800 31136
rect 79200 30880 80800 31000
rect -800 30608 800 30728
rect -800 30200 800 30320
rect 79200 30200 80800 30320
rect -800 29792 800 29912
rect -800 29384 800 29504
rect 79200 29520 80800 29640
rect -800 28976 800 29096
rect 79200 28976 80800 29096
rect -800 28568 800 28688
rect -800 28160 800 28280
rect 79200 28296 80800 28416
rect -800 27752 800 27872
rect 79200 27752 80800 27872
rect -800 27344 800 27464
rect -800 26936 800 27056
rect 79200 27072 80800 27192
rect -800 26664 800 26784
rect -800 26256 800 26376
rect 79200 26392 80800 26512
rect -800 25848 800 25968
rect 79200 25848 80800 25968
rect -800 25440 800 25560
rect -800 25032 800 25152
rect 79200 25168 80800 25288
rect -800 24624 800 24744
rect 79200 24624 80800 24744
rect -800 24216 800 24336
rect -800 23808 800 23928
rect 79200 23944 80800 24064
rect -800 23400 800 23520
rect 79200 23264 80800 23384
rect -800 22992 800 23112
rect -800 22584 800 22704
rect 79200 22720 80800 22840
rect -800 22176 800 22296
rect 79200 22040 80800 22160
rect -800 21768 800 21888
rect -800 21360 800 21480
rect 79200 21496 80800 21616
rect -800 20952 800 21072
rect 79200 20816 80800 20936
rect -800 20544 800 20664
rect -800 20136 800 20256
rect 79200 20272 80800 20392
rect -800 19728 800 19848
rect 79200 19592 80800 19712
rect -800 19320 800 19440
rect -800 18912 800 19032
rect 79200 18912 80800 19032
rect -800 18504 800 18624
rect 79200 18368 80800 18488
rect -800 18096 800 18216
rect -800 17824 800 17944
rect 79200 17688 80800 17808
rect -800 17416 800 17536
rect -800 17008 800 17128
rect 79200 17144 80800 17264
rect -800 16600 800 16720
rect 79200 16464 80800 16584
rect -800 16192 800 16312
rect -800 15784 800 15904
rect 79200 15784 80800 15904
rect -800 15376 800 15496
rect 79200 15240 80800 15360
rect -800 14968 800 15088
rect -800 14560 800 14680
rect 79200 14560 80800 14680
rect -800 14152 800 14272
rect 79200 14016 80800 14136
rect -800 13744 800 13864
rect -800 13336 800 13456
rect 79200 13336 80800 13456
rect -800 12928 800 13048
rect -800 12520 800 12640
rect 79200 12656 80800 12776
rect -800 12112 800 12232
rect 79200 12112 80800 12232
rect -800 11704 800 11824
rect -800 11296 800 11416
rect 79200 11432 80800 11552
rect -800 10888 800 11008
rect 79200 10888 80800 11008
rect -800 10480 800 10600
rect -800 10072 800 10192
rect 79200 10208 80800 10328
rect -800 9664 800 9784
rect 79200 9528 80800 9648
rect -800 9256 800 9376
rect -800 8984 800 9104
rect 79200 8984 80800 9104
rect -800 8576 800 8696
rect -800 8168 800 8288
rect 79200 8304 80800 8424
rect -800 7760 800 7880
rect 79200 7760 80800 7880
rect -800 7352 800 7472
rect -800 6944 800 7064
rect 79200 7080 80800 7200
rect -800 6536 800 6656
rect 79200 6400 80800 6520
rect -800 6128 800 6248
rect -800 5720 800 5840
rect 79200 5856 80800 5976
rect -800 5312 800 5432
rect 79200 5176 80800 5296
rect -800 4904 800 5024
rect -800 4496 800 4616
rect 79200 4632 80800 4752
rect -800 4088 800 4208
rect 79200 3952 80800 4072
rect -800 3680 800 3800
rect -800 3272 800 3392
rect 79200 3272 80800 3392
rect -800 2864 800 2984
rect 79200 2728 80800 2848
rect -800 2456 800 2576
rect -800 2048 800 2168
rect 79200 2048 80800 2168
rect -800 1640 800 1760
rect 79200 1504 80800 1624
rect -800 1232 800 1352
rect -800 824 800 944
rect 79200 824 80800 944
rect -800 416 800 536
rect 79200 280 80800 400
rect -800 144 800 264
<< obsm3 >>
rect 880 79768 79200 79797
rect 880 79624 79120 79768
rect 800 79496 79120 79624
rect 880 79488 79120 79496
rect 880 79216 79200 79488
rect 800 79088 79200 79216
rect 880 78808 79120 79088
rect 800 78680 79200 78808
rect 880 78544 79200 78680
rect 880 78400 79120 78544
rect 800 78272 79120 78400
rect 880 78264 79120 78272
rect 880 77992 79200 78264
rect 800 77864 79200 77992
rect 880 77584 79120 77864
rect 800 77456 79200 77584
rect 880 77320 79200 77456
rect 880 77176 79120 77320
rect 800 77048 79120 77176
rect 880 77040 79120 77048
rect 880 76768 79200 77040
rect 800 76640 79200 76768
rect 880 76360 79120 76640
rect 800 76232 79200 76360
rect 880 75960 79200 76232
rect 880 75952 79120 75960
rect 800 75824 79120 75952
rect 880 75680 79120 75824
rect 880 75544 79200 75680
rect 800 75416 79200 75544
rect 880 75136 79120 75416
rect 800 75008 79200 75136
rect 880 74736 79200 75008
rect 880 74728 79120 74736
rect 800 74600 79120 74728
rect 880 74456 79120 74600
rect 880 74320 79200 74456
rect 800 74192 79200 74320
rect 880 73912 79120 74192
rect 800 73784 79200 73912
rect 880 73512 79200 73784
rect 880 73504 79120 73512
rect 800 73376 79120 73504
rect 880 73232 79120 73376
rect 880 73096 79200 73232
rect 800 72968 79200 73096
rect 880 72832 79200 72968
rect 880 72688 79120 72832
rect 800 72560 79120 72688
rect 880 72552 79120 72560
rect 880 72288 79200 72552
rect 880 72280 79120 72288
rect 800 72152 79120 72280
rect 880 72008 79120 72152
rect 880 71872 79200 72008
rect 800 71744 79200 71872
rect 880 71608 79200 71744
rect 880 71464 79120 71608
rect 800 71336 79120 71464
rect 880 71328 79120 71336
rect 880 71064 79200 71328
rect 880 70784 79120 71064
rect 800 70656 79200 70784
rect 880 70384 79200 70656
rect 880 70376 79120 70384
rect 800 70248 79120 70376
rect 880 70104 79120 70248
rect 880 69968 79200 70104
rect 800 69840 79200 69968
rect 880 69704 79200 69840
rect 880 69560 79120 69704
rect 800 69432 79120 69560
rect 880 69424 79120 69432
rect 880 69160 79200 69424
rect 880 69152 79120 69160
rect 800 69024 79120 69152
rect 880 68880 79120 69024
rect 880 68744 79200 68880
rect 800 68616 79200 68744
rect 880 68480 79200 68616
rect 880 68336 79120 68480
rect 800 68208 79120 68336
rect 880 68200 79120 68208
rect 880 67936 79200 68200
rect 880 67928 79120 67936
rect 800 67800 79120 67928
rect 880 67656 79120 67800
rect 880 67520 79200 67656
rect 800 67392 79200 67520
rect 880 67256 79200 67392
rect 880 67112 79120 67256
rect 800 66984 79120 67112
rect 880 66976 79120 66984
rect 880 66704 79200 66976
rect 800 66576 79200 66704
rect 880 66296 79120 66576
rect 800 66168 79200 66296
rect 880 66032 79200 66168
rect 880 65888 79120 66032
rect 800 65760 79120 65888
rect 880 65752 79120 65760
rect 880 65480 79200 65752
rect 800 65352 79200 65480
rect 880 65072 79120 65352
rect 800 64944 79200 65072
rect 880 64808 79200 64944
rect 880 64664 79120 64808
rect 800 64536 79120 64664
rect 880 64528 79120 64536
rect 880 64256 79200 64528
rect 800 64128 79200 64256
rect 880 63848 79120 64128
rect 800 63720 79200 63848
rect 880 63448 79200 63720
rect 880 63440 79120 63448
rect 800 63312 79120 63440
rect 880 63168 79120 63312
rect 880 63032 79200 63168
rect 800 62904 79200 63032
rect 880 62624 79120 62904
rect 800 62496 79200 62624
rect 880 62224 79200 62496
rect 880 61944 79120 62224
rect 800 61816 79200 61944
rect 880 61680 79200 61816
rect 880 61536 79120 61680
rect 800 61408 79120 61536
rect 880 61400 79120 61408
rect 880 61128 79200 61400
rect 800 61000 79200 61128
rect 880 60720 79120 61000
rect 800 60592 79200 60720
rect 880 60456 79200 60592
rect 880 60312 79120 60456
rect 800 60184 79120 60312
rect 880 60176 79120 60184
rect 880 59904 79200 60176
rect 800 59776 79200 59904
rect 880 59496 79120 59776
rect 800 59368 79200 59496
rect 880 59096 79200 59368
rect 880 59088 79120 59096
rect 800 58960 79120 59088
rect 880 58816 79120 58960
rect 880 58680 79200 58816
rect 800 58552 79200 58680
rect 880 58272 79120 58552
rect 800 58144 79200 58272
rect 880 57872 79200 58144
rect 880 57864 79120 57872
rect 800 57736 79120 57864
rect 880 57592 79120 57736
rect 880 57456 79200 57592
rect 800 57328 79200 57456
rect 880 57048 79120 57328
rect 800 56920 79200 57048
rect 880 56648 79200 56920
rect 880 56640 79120 56648
rect 800 56512 79120 56640
rect 880 56368 79120 56512
rect 880 56232 79200 56368
rect 800 56104 79200 56232
rect 880 55968 79200 56104
rect 880 55824 79120 55968
rect 800 55696 79120 55824
rect 880 55688 79120 55696
rect 880 55424 79200 55688
rect 880 55416 79120 55424
rect 800 55288 79120 55416
rect 880 55144 79120 55288
rect 880 55008 79200 55144
rect 800 54880 79200 55008
rect 880 54744 79200 54880
rect 880 54600 79120 54744
rect 800 54472 79120 54600
rect 880 54464 79120 54472
rect 880 54200 79200 54464
rect 880 54192 79120 54200
rect 800 54064 79120 54192
rect 880 53920 79120 54064
rect 880 53784 79200 53920
rect 800 53656 79200 53784
rect 880 53520 79200 53656
rect 880 53240 79120 53520
rect 880 53104 79200 53240
rect 800 52976 79200 53104
rect 880 52840 79200 52976
rect 880 52696 79120 52840
rect 800 52568 79120 52696
rect 880 52560 79120 52568
rect 880 52296 79200 52560
rect 880 52288 79120 52296
rect 800 52160 79120 52288
rect 880 52016 79120 52160
rect 880 51880 79200 52016
rect 800 51752 79200 51880
rect 880 51616 79200 51752
rect 880 51472 79120 51616
rect 800 51344 79120 51472
rect 880 51336 79120 51344
rect 880 51072 79200 51336
rect 880 51064 79120 51072
rect 800 50936 79120 51064
rect 880 50792 79120 50936
rect 880 50656 79200 50792
rect 800 50528 79200 50656
rect 880 50392 79200 50528
rect 880 50248 79120 50392
rect 800 50120 79120 50248
rect 880 50112 79120 50120
rect 880 49840 79200 50112
rect 800 49712 79200 49840
rect 880 49432 79120 49712
rect 800 49304 79200 49432
rect 880 49168 79200 49304
rect 880 49024 79120 49168
rect 800 48896 79120 49024
rect 880 48888 79120 48896
rect 880 48616 79200 48888
rect 800 48488 79200 48616
rect 880 48208 79120 48488
rect 800 48080 79200 48208
rect 880 47944 79200 48080
rect 880 47800 79120 47944
rect 800 47672 79120 47800
rect 880 47664 79120 47672
rect 880 47392 79200 47664
rect 800 47264 79200 47392
rect 880 46984 79120 47264
rect 800 46856 79200 46984
rect 880 46584 79200 46856
rect 880 46576 79120 46584
rect 800 46448 79120 46576
rect 880 46304 79120 46448
rect 880 46168 79200 46304
rect 800 46040 79200 46168
rect 880 45760 79120 46040
rect 800 45632 79200 45760
rect 880 45360 79200 45632
rect 880 45352 79120 45360
rect 800 45224 79120 45352
rect 880 45080 79120 45224
rect 880 44944 79200 45080
rect 800 44816 79200 44944
rect 880 44536 79120 44816
rect 880 44264 79200 44536
rect 800 44136 79200 44264
rect 880 43856 79120 44136
rect 800 43728 79200 43856
rect 880 43456 79200 43728
rect 880 43448 79120 43456
rect 800 43320 79120 43448
rect 880 43176 79120 43320
rect 880 43040 79200 43176
rect 800 42912 79200 43040
rect 880 42632 79120 42912
rect 800 42504 79200 42632
rect 880 42232 79200 42504
rect 880 42224 79120 42232
rect 800 42096 79120 42224
rect 880 41952 79120 42096
rect 880 41816 79200 41952
rect 800 41688 79200 41816
rect 880 41408 79120 41688
rect 800 41280 79200 41408
rect 880 41008 79200 41280
rect 880 41000 79120 41008
rect 800 40872 79120 41000
rect 880 40728 79120 40872
rect 880 40592 79200 40728
rect 800 40464 79200 40592
rect 880 40184 79120 40464
rect 800 40056 79200 40184
rect 880 39784 79200 40056
rect 880 39776 79120 39784
rect 800 39648 79120 39776
rect 880 39504 79120 39648
rect 880 39368 79200 39504
rect 800 39240 79200 39368
rect 880 39104 79200 39240
rect 880 38960 79120 39104
rect 800 38832 79120 38960
rect 880 38824 79120 38832
rect 880 38560 79200 38824
rect 880 38552 79120 38560
rect 800 38424 79120 38552
rect 880 38280 79120 38424
rect 880 38144 79200 38280
rect 800 38016 79200 38144
rect 880 37880 79200 38016
rect 880 37736 79120 37880
rect 800 37608 79120 37736
rect 880 37600 79120 37608
rect 880 37336 79200 37600
rect 880 37328 79120 37336
rect 800 37200 79120 37328
rect 880 37056 79120 37200
rect 880 36920 79200 37056
rect 800 36792 79200 36920
rect 880 36656 79200 36792
rect 880 36512 79120 36656
rect 800 36384 79120 36512
rect 880 36376 79120 36384
rect 880 36104 79200 36376
rect 800 35976 79200 36104
rect 880 35696 79120 35976
rect 880 35432 79200 35696
rect 880 35424 79120 35432
rect 800 35296 79120 35424
rect 880 35152 79120 35296
rect 880 35016 79200 35152
rect 800 34888 79200 35016
rect 880 34752 79200 34888
rect 880 34608 79120 34752
rect 800 34480 79120 34608
rect 880 34472 79120 34480
rect 880 34208 79200 34472
rect 880 34200 79120 34208
rect 800 34072 79120 34200
rect 880 33928 79120 34072
rect 880 33792 79200 33928
rect 800 33664 79200 33792
rect 880 33528 79200 33664
rect 880 33384 79120 33528
rect 800 33256 79120 33384
rect 880 33248 79120 33256
rect 880 32976 79200 33248
rect 800 32848 79200 32976
rect 880 32568 79120 32848
rect 800 32440 79200 32568
rect 880 32304 79200 32440
rect 880 32160 79120 32304
rect 800 32032 79120 32160
rect 880 32024 79120 32032
rect 880 31752 79200 32024
rect 800 31624 79200 31752
rect 880 31344 79120 31624
rect 800 31216 79200 31344
rect 880 31080 79200 31216
rect 880 30936 79120 31080
rect 800 30808 79120 30936
rect 880 30800 79120 30808
rect 880 30528 79200 30800
rect 800 30400 79200 30528
rect 880 30120 79120 30400
rect 800 29992 79200 30120
rect 880 29720 79200 29992
rect 880 29712 79120 29720
rect 800 29584 79120 29712
rect 880 29440 79120 29584
rect 880 29304 79200 29440
rect 800 29176 79200 29304
rect 880 28896 79120 29176
rect 800 28768 79200 28896
rect 880 28496 79200 28768
rect 880 28488 79120 28496
rect 800 28360 79120 28488
rect 880 28216 79120 28360
rect 880 28080 79200 28216
rect 800 27952 79200 28080
rect 880 27672 79120 27952
rect 800 27544 79200 27672
rect 880 27272 79200 27544
rect 880 27264 79120 27272
rect 800 27136 79120 27264
rect 880 26992 79120 27136
rect 880 26592 79200 26992
rect 880 26584 79120 26592
rect 800 26456 79120 26584
rect 880 26312 79120 26456
rect 880 26176 79200 26312
rect 800 26048 79200 26176
rect 880 25768 79120 26048
rect 800 25640 79200 25768
rect 880 25368 79200 25640
rect 880 25360 79120 25368
rect 800 25232 79120 25360
rect 880 25088 79120 25232
rect 880 24952 79200 25088
rect 800 24824 79200 24952
rect 880 24544 79120 24824
rect 800 24416 79200 24544
rect 880 24144 79200 24416
rect 880 24136 79120 24144
rect 800 24008 79120 24136
rect 880 23864 79120 24008
rect 880 23728 79200 23864
rect 800 23600 79200 23728
rect 880 23464 79200 23600
rect 880 23320 79120 23464
rect 800 23192 79120 23320
rect 880 23184 79120 23192
rect 880 22920 79200 23184
rect 880 22912 79120 22920
rect 800 22784 79120 22912
rect 880 22640 79120 22784
rect 880 22504 79200 22640
rect 800 22376 79200 22504
rect 880 22240 79200 22376
rect 880 22096 79120 22240
rect 800 21968 79120 22096
rect 880 21960 79120 21968
rect 880 21696 79200 21960
rect 880 21688 79120 21696
rect 800 21560 79120 21688
rect 880 21416 79120 21560
rect 880 21280 79200 21416
rect 800 21152 79200 21280
rect 880 21016 79200 21152
rect 880 20872 79120 21016
rect 800 20744 79120 20872
rect 880 20736 79120 20744
rect 880 20472 79200 20736
rect 880 20464 79120 20472
rect 800 20336 79120 20464
rect 880 20192 79120 20336
rect 880 20056 79200 20192
rect 800 19928 79200 20056
rect 880 19792 79200 19928
rect 880 19648 79120 19792
rect 800 19520 79120 19648
rect 880 19512 79120 19520
rect 880 19240 79200 19512
rect 800 19112 79200 19240
rect 880 18832 79120 19112
rect 800 18704 79200 18832
rect 880 18568 79200 18704
rect 880 18424 79120 18568
rect 800 18296 79120 18424
rect 880 18288 79120 18296
rect 880 17888 79200 18288
rect 880 17744 79120 17888
rect 800 17616 79120 17744
rect 880 17608 79120 17616
rect 880 17344 79200 17608
rect 880 17336 79120 17344
rect 800 17208 79120 17336
rect 880 17064 79120 17208
rect 880 16928 79200 17064
rect 800 16800 79200 16928
rect 880 16664 79200 16800
rect 880 16520 79120 16664
rect 800 16392 79120 16520
rect 880 16384 79120 16392
rect 880 16112 79200 16384
rect 800 15984 79200 16112
rect 880 15704 79120 15984
rect 800 15576 79200 15704
rect 880 15440 79200 15576
rect 880 15296 79120 15440
rect 800 15168 79120 15296
rect 880 15160 79120 15168
rect 880 14888 79200 15160
rect 800 14760 79200 14888
rect 880 14480 79120 14760
rect 800 14352 79200 14480
rect 880 14216 79200 14352
rect 880 14072 79120 14216
rect 800 13944 79120 14072
rect 880 13936 79120 13944
rect 880 13664 79200 13936
rect 800 13536 79200 13664
rect 880 13256 79120 13536
rect 800 13128 79200 13256
rect 880 12856 79200 13128
rect 880 12848 79120 12856
rect 800 12720 79120 12848
rect 880 12576 79120 12720
rect 880 12440 79200 12576
rect 800 12312 79200 12440
rect 880 12032 79120 12312
rect 800 11904 79200 12032
rect 880 11632 79200 11904
rect 880 11624 79120 11632
rect 800 11496 79120 11624
rect 880 11352 79120 11496
rect 880 11216 79200 11352
rect 800 11088 79200 11216
rect 880 10808 79120 11088
rect 800 10680 79200 10808
rect 880 10408 79200 10680
rect 880 10400 79120 10408
rect 800 10272 79120 10400
rect 880 10128 79120 10272
rect 880 9992 79200 10128
rect 800 9864 79200 9992
rect 880 9728 79200 9864
rect 880 9584 79120 9728
rect 800 9456 79120 9584
rect 880 9448 79120 9456
rect 880 9184 79200 9448
rect 880 8904 79120 9184
rect 800 8776 79200 8904
rect 880 8504 79200 8776
rect 880 8496 79120 8504
rect 800 8368 79120 8496
rect 880 8224 79120 8368
rect 880 8088 79200 8224
rect 800 7960 79200 8088
rect 880 7680 79120 7960
rect 800 7552 79200 7680
rect 880 7280 79200 7552
rect 880 7272 79120 7280
rect 800 7144 79120 7272
rect 880 7000 79120 7144
rect 880 6864 79200 7000
rect 800 6736 79200 6864
rect 880 6600 79200 6736
rect 880 6456 79120 6600
rect 800 6328 79120 6456
rect 880 6320 79120 6328
rect 880 6056 79200 6320
rect 880 6048 79120 6056
rect 800 5920 79120 6048
rect 880 5776 79120 5920
rect 880 5640 79200 5776
rect 800 5512 79200 5640
rect 880 5376 79200 5512
rect 880 5232 79120 5376
rect 800 5104 79120 5232
rect 880 5096 79120 5104
rect 880 4832 79200 5096
rect 880 4824 79120 4832
rect 800 4696 79120 4824
rect 880 4552 79120 4696
rect 880 4416 79200 4552
rect 800 4288 79200 4416
rect 880 4152 79200 4288
rect 880 4008 79120 4152
rect 800 3880 79120 4008
rect 880 3872 79120 3880
rect 880 3600 79200 3872
rect 800 3472 79200 3600
rect 880 3192 79120 3472
rect 800 3064 79200 3192
rect 880 2928 79200 3064
rect 880 2784 79120 2928
rect 800 2656 79120 2784
rect 880 2648 79120 2656
rect 880 2376 79200 2648
rect 800 2248 79200 2376
rect 880 1968 79120 2248
rect 800 1840 79200 1968
rect 880 1704 79200 1840
rect 880 1560 79120 1704
rect 800 1432 79120 1560
rect 880 1424 79120 1432
rect 880 1152 79200 1424
rect 800 1024 79200 1152
rect 880 744 79120 1024
rect 800 616 79200 744
rect 880 480 79200 616
rect 880 307 79120 480
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< labels >>
rlabel metal2 s 110 79200 166 80800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 3330 79200 3386 80800 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 3698 79200 3754 80800 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 3974 79200 4030 80800 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 4342 79200 4398 80800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 4710 79200 4766 80800 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 4986 79200 5042 80800 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 5354 79200 5410 80800 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 5630 79200 5686 80800 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 5998 79200 6054 80800 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 6366 79200 6422 80800 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 386 79200 442 80800 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 6642 79200 6698 80800 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 7010 79200 7066 80800 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 7286 79200 7342 80800 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 7654 79200 7710 80800 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 7930 79200 7986 80800 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 8298 79200 8354 80800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 8666 79200 8722 80800 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 8942 79200 8998 80800 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 9310 79200 9366 80800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 9586 79200 9642 80800 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 754 79200 810 80800 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 9954 79200 10010 80800 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 10230 79200 10286 80800 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 10598 79200 10654 80800 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 10966 79200 11022 80800 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 11242 79200 11298 80800 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 11610 79200 11666 80800 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 11886 79200 11942 80800 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 12254 79200 12310 80800 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 1030 79200 1086 80800 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 1398 79200 1454 80800 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 1674 79200 1730 80800 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 2042 79200 2098 80800 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 2410 79200 2466 80800 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 2686 79200 2742 80800 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 3054 79200 3110 80800 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 25134 79200 25190 80800 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 28354 79200 28410 80800 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 28722 79200 28778 80800 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 29090 79200 29146 80800 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 29366 79200 29422 80800 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 29734 79200 29790 80800 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 30010 79200 30066 80800 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 30378 79200 30434 80800 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 30654 79200 30710 80800 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 31022 79200 31078 80800 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 31390 79200 31446 80800 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 25410 79200 25466 80800 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 31666 79200 31722 80800 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 32034 79200 32090 80800 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 32310 79200 32366 80800 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 32678 79200 32734 80800 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 33046 79200 33102 80800 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 33322 79200 33378 80800 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 33690 79200 33746 80800 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 33966 79200 34022 80800 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 34334 79200 34390 80800 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 34610 79200 34666 80800 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 25778 79200 25834 80800 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 34978 79200 35034 80800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 35346 79200 35402 80800 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 35622 79200 35678 80800 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 35990 79200 36046 80800 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 36266 79200 36322 80800 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 36634 79200 36690 80800 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 36910 79200 36966 80800 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 37278 79200 37334 80800 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 26054 79200 26110 80800 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 26422 79200 26478 80800 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 26790 79200 26846 80800 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 27066 79200 27122 80800 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 27434 79200 27490 80800 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 27710 79200 27766 80800 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 28078 79200 28134 80800 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 12622 79200 12678 80800 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 15842 79200 15898 80800 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 16210 79200 16266 80800 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 16578 79200 16634 80800 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 16854 79200 16910 80800 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 17222 79200 17278 80800 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 17498 79200 17554 80800 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 17866 79200 17922 80800 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 18142 79200 18198 80800 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 18510 79200 18566 80800 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 18878 79200 18934 80800 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 12898 79200 12954 80800 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 19154 79200 19210 80800 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 19522 79200 19578 80800 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 19798 79200 19854 80800 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 20166 79200 20222 80800 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 20442 79200 20498 80800 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 20810 79200 20866 80800 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 21178 79200 21234 80800 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 21454 79200 21510 80800 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 21822 79200 21878 80800 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 22098 79200 22154 80800 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 13266 79200 13322 80800 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 22466 79200 22522 80800 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 22834 79200 22890 80800 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 23110 79200 23166 80800 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 23478 79200 23534 80800 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 23754 79200 23810 80800 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 24122 79200 24178 80800 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 24398 79200 24454 80800 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 24766 79200 24822 80800 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 13542 79200 13598 80800 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 13910 79200 13966 80800 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14186 79200 14242 80800 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 14554 79200 14610 80800 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 14922 79200 14978 80800 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 15198 79200 15254 80800 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 15566 79200 15622 80800 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s -800 27344 800 27464 4 irq[0]
port 115 nsew signal output
rlabel metal3 s -800 27752 800 27872 4 irq[1]
port 116 nsew signal output
rlabel metal3 s -800 28160 800 28280 4 irq[2]
port 117 nsew signal output
rlabel metal2 s 294 -800 350 800 8 la_data_out[0]
port 118 nsew signal output
rlabel metal2 s 62762 -800 62818 800 8 la_data_out[100]
port 119 nsew signal output
rlabel metal2 s 63406 -800 63462 800 8 la_data_out[101]
port 120 nsew signal output
rlabel metal2 s 64050 -800 64106 800 8 la_data_out[102]
port 121 nsew signal output
rlabel metal2 s 64694 -800 64750 800 8 la_data_out[103]
port 122 nsew signal output
rlabel metal2 s 65246 -800 65302 800 8 la_data_out[104]
port 123 nsew signal output
rlabel metal2 s 65890 -800 65946 800 8 la_data_out[105]
port 124 nsew signal output
rlabel metal2 s 66534 -800 66590 800 8 la_data_out[106]
port 125 nsew signal output
rlabel metal2 s 67178 -800 67234 800 8 la_data_out[107]
port 126 nsew signal output
rlabel metal2 s 67822 -800 67878 800 8 la_data_out[108]
port 127 nsew signal output
rlabel metal2 s 68374 -800 68430 800 8 la_data_out[109]
port 128 nsew signal output
rlabel metal2 s 6458 -800 6514 800 8 la_data_out[10]
port 129 nsew signal output
rlabel metal2 s 69018 -800 69074 800 8 la_data_out[110]
port 130 nsew signal output
rlabel metal2 s 69662 -800 69718 800 8 la_data_out[111]
port 131 nsew signal output
rlabel metal2 s 70306 -800 70362 800 8 la_data_out[112]
port 132 nsew signal output
rlabel metal2 s 70950 -800 71006 800 8 la_data_out[113]
port 133 nsew signal output
rlabel metal2 s 71502 -800 71558 800 8 la_data_out[114]
port 134 nsew signal output
rlabel metal2 s 72146 -800 72202 800 8 la_data_out[115]
port 135 nsew signal output
rlabel metal2 s 72790 -800 72846 800 8 la_data_out[116]
port 136 nsew signal output
rlabel metal2 s 73434 -800 73490 800 8 la_data_out[117]
port 137 nsew signal output
rlabel metal2 s 74078 -800 74134 800 8 la_data_out[118]
port 138 nsew signal output
rlabel metal2 s 74630 -800 74686 800 8 la_data_out[119]
port 139 nsew signal output
rlabel metal2 s 7102 -800 7158 800 8 la_data_out[11]
port 140 nsew signal output
rlabel metal2 s 75274 -800 75330 800 8 la_data_out[120]
port 141 nsew signal output
rlabel metal2 s 75918 -800 75974 800 8 la_data_out[121]
port 142 nsew signal output
rlabel metal2 s 76562 -800 76618 800 8 la_data_out[122]
port 143 nsew signal output
rlabel metal2 s 77206 -800 77262 800 8 la_data_out[123]
port 144 nsew signal output
rlabel metal2 s 77758 -800 77814 800 8 la_data_out[124]
port 145 nsew signal output
rlabel metal2 s 78402 -800 78458 800 8 la_data_out[125]
port 146 nsew signal output
rlabel metal2 s 79046 -800 79102 800 8 la_data_out[126]
port 147 nsew signal output
rlabel metal2 s 79690 -800 79746 800 8 la_data_out[127]
port 148 nsew signal output
rlabel metal2 s 7746 -800 7802 800 8 la_data_out[12]
port 149 nsew signal output
rlabel metal2 s 8390 -800 8446 800 8 la_data_out[13]
port 150 nsew signal output
rlabel metal2 s 9034 -800 9090 800 8 la_data_out[14]
port 151 nsew signal output
rlabel metal2 s 9586 -800 9642 800 8 la_data_out[15]
port 152 nsew signal output
rlabel metal2 s 10230 -800 10286 800 8 la_data_out[16]
port 153 nsew signal output
rlabel metal2 s 10874 -800 10930 800 8 la_data_out[17]
port 154 nsew signal output
rlabel metal2 s 11518 -800 11574 800 8 la_data_out[18]
port 155 nsew signal output
rlabel metal2 s 12162 -800 12218 800 8 la_data_out[19]
port 156 nsew signal output
rlabel metal2 s 846 -800 902 800 8 la_data_out[1]
port 157 nsew signal output
rlabel metal2 s 12714 -800 12770 800 8 la_data_out[20]
port 158 nsew signal output
rlabel metal2 s 13358 -800 13414 800 8 la_data_out[21]
port 159 nsew signal output
rlabel metal2 s 14002 -800 14058 800 8 la_data_out[22]
port 160 nsew signal output
rlabel metal2 s 14646 -800 14702 800 8 la_data_out[23]
port 161 nsew signal output
rlabel metal2 s 15290 -800 15346 800 8 la_data_out[24]
port 162 nsew signal output
rlabel metal2 s 15842 -800 15898 800 8 la_data_out[25]
port 163 nsew signal output
rlabel metal2 s 16486 -800 16542 800 8 la_data_out[26]
port 164 nsew signal output
rlabel metal2 s 17130 -800 17186 800 8 la_data_out[27]
port 165 nsew signal output
rlabel metal2 s 17774 -800 17830 800 8 la_data_out[28]
port 166 nsew signal output
rlabel metal2 s 18418 -800 18474 800 8 la_data_out[29]
port 167 nsew signal output
rlabel metal2 s 1490 -800 1546 800 8 la_data_out[2]
port 168 nsew signal output
rlabel metal2 s 18970 -800 19026 800 8 la_data_out[30]
port 169 nsew signal output
rlabel metal2 s 19614 -800 19670 800 8 la_data_out[31]
port 170 nsew signal output
rlabel metal2 s 20258 -800 20314 800 8 la_data_out[32]
port 171 nsew signal output
rlabel metal2 s 20902 -800 20958 800 8 la_data_out[33]
port 172 nsew signal output
rlabel metal2 s 21546 -800 21602 800 8 la_data_out[34]
port 173 nsew signal output
rlabel metal2 s 22098 -800 22154 800 8 la_data_out[35]
port 174 nsew signal output
rlabel metal2 s 22742 -800 22798 800 8 la_data_out[36]
port 175 nsew signal output
rlabel metal2 s 23386 -800 23442 800 8 la_data_out[37]
port 176 nsew signal output
rlabel metal2 s 24030 -800 24086 800 8 la_data_out[38]
port 177 nsew signal output
rlabel metal2 s 24674 -800 24730 800 8 la_data_out[39]
port 178 nsew signal output
rlabel metal2 s 2134 -800 2190 800 8 la_data_out[3]
port 179 nsew signal output
rlabel metal2 s 25226 -800 25282 800 8 la_data_out[40]
port 180 nsew signal output
rlabel metal2 s 25870 -800 25926 800 8 la_data_out[41]
port 181 nsew signal output
rlabel metal2 s 26514 -800 26570 800 8 la_data_out[42]
port 182 nsew signal output
rlabel metal2 s 27158 -800 27214 800 8 la_data_out[43]
port 183 nsew signal output
rlabel metal2 s 27802 -800 27858 800 8 la_data_out[44]
port 184 nsew signal output
rlabel metal2 s 28354 -800 28410 800 8 la_data_out[45]
port 185 nsew signal output
rlabel metal2 s 28998 -800 29054 800 8 la_data_out[46]
port 186 nsew signal output
rlabel metal2 s 29642 -800 29698 800 8 la_data_out[47]
port 187 nsew signal output
rlabel metal2 s 30286 -800 30342 800 8 la_data_out[48]
port 188 nsew signal output
rlabel metal2 s 30930 -800 30986 800 8 la_data_out[49]
port 189 nsew signal output
rlabel metal2 s 2778 -800 2834 800 8 la_data_out[4]
port 190 nsew signal output
rlabel metal2 s 31482 -800 31538 800 8 la_data_out[50]
port 191 nsew signal output
rlabel metal2 s 32126 -800 32182 800 8 la_data_out[51]
port 192 nsew signal output
rlabel metal2 s 32770 -800 32826 800 8 la_data_out[52]
port 193 nsew signal output
rlabel metal2 s 33414 -800 33470 800 8 la_data_out[53]
port 194 nsew signal output
rlabel metal2 s 34058 -800 34114 800 8 la_data_out[54]
port 195 nsew signal output
rlabel metal2 s 34610 -800 34666 800 8 la_data_out[55]
port 196 nsew signal output
rlabel metal2 s 35254 -800 35310 800 8 la_data_out[56]
port 197 nsew signal output
rlabel metal2 s 35898 -800 35954 800 8 la_data_out[57]
port 198 nsew signal output
rlabel metal2 s 36542 -800 36598 800 8 la_data_out[58]
port 199 nsew signal output
rlabel metal2 s 37186 -800 37242 800 8 la_data_out[59]
port 200 nsew signal output
rlabel metal2 s 3330 -800 3386 800 8 la_data_out[5]
port 201 nsew signal output
rlabel metal2 s 37738 -800 37794 800 8 la_data_out[60]
port 202 nsew signal output
rlabel metal2 s 38382 -800 38438 800 8 la_data_out[61]
port 203 nsew signal output
rlabel metal2 s 39026 -800 39082 800 8 la_data_out[62]
port 204 nsew signal output
rlabel metal2 s 39670 -800 39726 800 8 la_data_out[63]
port 205 nsew signal output
rlabel metal2 s 40314 -800 40370 800 8 la_data_out[64]
port 206 nsew signal output
rlabel metal2 s 40866 -800 40922 800 8 la_data_out[65]
port 207 nsew signal output
rlabel metal2 s 41510 -800 41566 800 8 la_data_out[66]
port 208 nsew signal output
rlabel metal2 s 42154 -800 42210 800 8 la_data_out[67]
port 209 nsew signal output
rlabel metal2 s 42798 -800 42854 800 8 la_data_out[68]
port 210 nsew signal output
rlabel metal2 s 43350 -800 43406 800 8 la_data_out[69]
port 211 nsew signal output
rlabel metal2 s 3974 -800 4030 800 8 la_data_out[6]
port 212 nsew signal output
rlabel metal2 s 43994 -800 44050 800 8 la_data_out[70]
port 213 nsew signal output
rlabel metal2 s 44638 -800 44694 800 8 la_data_out[71]
port 214 nsew signal output
rlabel metal2 s 45282 -800 45338 800 8 la_data_out[72]
port 215 nsew signal output
rlabel metal2 s 45926 -800 45982 800 8 la_data_out[73]
port 216 nsew signal output
rlabel metal2 s 46478 -800 46534 800 8 la_data_out[74]
port 217 nsew signal output
rlabel metal2 s 47122 -800 47178 800 8 la_data_out[75]
port 218 nsew signal output
rlabel metal2 s 47766 -800 47822 800 8 la_data_out[76]
port 219 nsew signal output
rlabel metal2 s 48410 -800 48466 800 8 la_data_out[77]
port 220 nsew signal output
rlabel metal2 s 49054 -800 49110 800 8 la_data_out[78]
port 221 nsew signal output
rlabel metal2 s 49606 -800 49662 800 8 la_data_out[79]
port 222 nsew signal output
rlabel metal2 s 4618 -800 4674 800 8 la_data_out[7]
port 223 nsew signal output
rlabel metal2 s 50250 -800 50306 800 8 la_data_out[80]
port 224 nsew signal output
rlabel metal2 s 50894 -800 50950 800 8 la_data_out[81]
port 225 nsew signal output
rlabel metal2 s 51538 -800 51594 800 8 la_data_out[82]
port 226 nsew signal output
rlabel metal2 s 52182 -800 52238 800 8 la_data_out[83]
port 227 nsew signal output
rlabel metal2 s 52734 -800 52790 800 8 la_data_out[84]
port 228 nsew signal output
rlabel metal2 s 53378 -800 53434 800 8 la_data_out[85]
port 229 nsew signal output
rlabel metal2 s 54022 -800 54078 800 8 la_data_out[86]
port 230 nsew signal output
rlabel metal2 s 54666 -800 54722 800 8 la_data_out[87]
port 231 nsew signal output
rlabel metal2 s 55310 -800 55366 800 8 la_data_out[88]
port 232 nsew signal output
rlabel metal2 s 55862 -800 55918 800 8 la_data_out[89]
port 233 nsew signal output
rlabel metal2 s 5262 -800 5318 800 8 la_data_out[8]
port 234 nsew signal output
rlabel metal2 s 56506 -800 56562 800 8 la_data_out[90]
port 235 nsew signal output
rlabel metal2 s 57150 -800 57206 800 8 la_data_out[91]
port 236 nsew signal output
rlabel metal2 s 57794 -800 57850 800 8 la_data_out[92]
port 237 nsew signal output
rlabel metal2 s 58438 -800 58494 800 8 la_data_out[93]
port 238 nsew signal output
rlabel metal2 s 58990 -800 59046 800 8 la_data_out[94]
port 239 nsew signal output
rlabel metal2 s 59634 -800 59690 800 8 la_data_out[95]
port 240 nsew signal output
rlabel metal2 s 60278 -800 60334 800 8 la_data_out[96]
port 241 nsew signal output
rlabel metal2 s 60922 -800 60978 800 8 la_data_out[97]
port 242 nsew signal output
rlabel metal2 s 61566 -800 61622 800 8 la_data_out[98]
port 243 nsew signal output
rlabel metal2 s 62118 -800 62174 800 8 la_data_out[99]
port 244 nsew signal output
rlabel metal2 s 5906 -800 5962 800 8 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 37646 79200 37702 80800 6 m_wb_rst_i[0]
port 246 nsew signal output
rlabel metal2 s 40866 79200 40922 80800 6 m_wb_rst_i[10]
port 247 nsew signal output
rlabel metal2 s 37922 79200 37978 80800 6 m_wb_rst_i[1]
port 248 nsew signal output
rlabel metal2 s 38290 79200 38346 80800 6 m_wb_rst_i[2]
port 249 nsew signal output
rlabel metal2 s 38566 79200 38622 80800 6 m_wb_rst_i[3]
port 250 nsew signal output
rlabel metal2 s 38934 79200 38990 80800 6 m_wb_rst_i[4]
port 251 nsew signal output
rlabel metal2 s 39302 79200 39358 80800 6 m_wb_rst_i[5]
port 252 nsew signal output
rlabel metal2 s 39578 79200 39634 80800 6 m_wb_rst_i[6]
port 253 nsew signal output
rlabel metal2 s 39946 79200 40002 80800 6 m_wb_rst_i[7]
port 254 nsew signal output
rlabel metal2 s 40222 79200 40278 80800 6 m_wb_rst_i[8]
port 255 nsew signal output
rlabel metal2 s 40590 79200 40646 80800 6 m_wb_rst_i[9]
port 256 nsew signal output
rlabel metal2 s 44822 79200 44878 80800 6 m_wbs_ack_o[0]
port 257 nsew signal input
rlabel metal2 s 48134 79200 48190 80800 6 m_wbs_ack_o[10]
port 258 nsew signal input
rlabel metal2 s 45190 79200 45246 80800 6 m_wbs_ack_o[1]
port 259 nsew signal input
rlabel metal2 s 45558 79200 45614 80800 6 m_wbs_ack_o[2]
port 260 nsew signal input
rlabel metal2 s 45834 79200 45890 80800 6 m_wbs_ack_o[3]
port 261 nsew signal input
rlabel metal2 s 46202 79200 46258 80800 6 m_wbs_ack_o[4]
port 262 nsew signal input
rlabel metal2 s 46478 79200 46534 80800 6 m_wbs_ack_o[5]
port 263 nsew signal input
rlabel metal2 s 46846 79200 46902 80800 6 m_wbs_ack_o[6]
port 264 nsew signal input
rlabel metal2 s 47122 79200 47178 80800 6 m_wbs_ack_o[7]
port 265 nsew signal input
rlabel metal2 s 47490 79200 47546 80800 6 m_wbs_ack_o[8]
port 266 nsew signal input
rlabel metal2 s 47858 79200 47914 80800 6 m_wbs_ack_o[9]
port 267 nsew signal input
rlabel metal3 s -800 28568 800 28688 4 m_wbs_dat_o_0[0]
port 268 nsew signal input
rlabel metal3 s -800 32648 800 32768 4 m_wbs_dat_o_0[10]
port 269 nsew signal input
rlabel metal3 s -800 33056 800 33176 4 m_wbs_dat_o_0[11]
port 270 nsew signal input
rlabel metal3 s -800 33464 800 33584 4 m_wbs_dat_o_0[12]
port 271 nsew signal input
rlabel metal3 s -800 33872 800 33992 4 m_wbs_dat_o_0[13]
port 272 nsew signal input
rlabel metal3 s -800 34280 800 34400 4 m_wbs_dat_o_0[14]
port 273 nsew signal input
rlabel metal3 s -800 34688 800 34808 4 m_wbs_dat_o_0[15]
port 274 nsew signal input
rlabel metal3 s -800 35096 800 35216 4 m_wbs_dat_o_0[16]
port 275 nsew signal input
rlabel metal3 s -800 35504 800 35624 4 m_wbs_dat_o_0[17]
port 276 nsew signal input
rlabel metal3 s -800 35776 800 35896 4 m_wbs_dat_o_0[18]
port 277 nsew signal input
rlabel metal3 s -800 36184 800 36304 4 m_wbs_dat_o_0[19]
port 278 nsew signal input
rlabel metal3 s -800 28976 800 29096 4 m_wbs_dat_o_0[1]
port 279 nsew signal input
rlabel metal3 s -800 36592 800 36712 4 m_wbs_dat_o_0[20]
port 280 nsew signal input
rlabel metal3 s -800 37000 800 37120 4 m_wbs_dat_o_0[21]
port 281 nsew signal input
rlabel metal3 s -800 37408 800 37528 4 m_wbs_dat_o_0[22]
port 282 nsew signal input
rlabel metal3 s -800 37816 800 37936 4 m_wbs_dat_o_0[23]
port 283 nsew signal input
rlabel metal3 s -800 38224 800 38344 4 m_wbs_dat_o_0[24]
port 284 nsew signal input
rlabel metal3 s -800 38632 800 38752 4 m_wbs_dat_o_0[25]
port 285 nsew signal input
rlabel metal3 s -800 39040 800 39160 4 m_wbs_dat_o_0[26]
port 286 nsew signal input
rlabel metal3 s -800 39448 800 39568 4 m_wbs_dat_o_0[27]
port 287 nsew signal input
rlabel metal3 s -800 39856 800 39976 4 m_wbs_dat_o_0[28]
port 288 nsew signal input
rlabel metal3 s -800 40264 800 40384 4 m_wbs_dat_o_0[29]
port 289 nsew signal input
rlabel metal3 s -800 29384 800 29504 4 m_wbs_dat_o_0[2]
port 290 nsew signal input
rlabel metal3 s -800 40672 800 40792 4 m_wbs_dat_o_0[30]
port 291 nsew signal input
rlabel metal3 s -800 41080 800 41200 4 m_wbs_dat_o_0[31]
port 292 nsew signal input
rlabel metal3 s -800 29792 800 29912 4 m_wbs_dat_o_0[3]
port 293 nsew signal input
rlabel metal3 s -800 30200 800 30320 4 m_wbs_dat_o_0[4]
port 294 nsew signal input
rlabel metal3 s -800 30608 800 30728 4 m_wbs_dat_o_0[5]
port 295 nsew signal input
rlabel metal3 s -800 31016 800 31136 4 m_wbs_dat_o_0[6]
port 296 nsew signal input
rlabel metal3 s -800 31424 800 31544 4 m_wbs_dat_o_0[7]
port 297 nsew signal input
rlabel metal3 s -800 31832 800 31952 4 m_wbs_dat_o_0[8]
port 298 nsew signal input
rlabel metal3 s -800 32240 800 32360 4 m_wbs_dat_o_0[9]
port 299 nsew signal input
rlabel metal3 s 79200 60256 80800 60376 6 m_wbs_dat_o_10[0]
port 300 nsew signal input
rlabel metal3 s 79200 66376 80800 66496 6 m_wbs_dat_o_10[10]
port 301 nsew signal input
rlabel metal3 s 79200 67056 80800 67176 6 m_wbs_dat_o_10[11]
port 302 nsew signal input
rlabel metal3 s 79200 67736 80800 67856 6 m_wbs_dat_o_10[12]
port 303 nsew signal input
rlabel metal3 s 79200 68280 80800 68400 6 m_wbs_dat_o_10[13]
port 304 nsew signal input
rlabel metal3 s 79200 68960 80800 69080 6 m_wbs_dat_o_10[14]
port 305 nsew signal input
rlabel metal3 s 79200 69504 80800 69624 6 m_wbs_dat_o_10[15]
port 306 nsew signal input
rlabel metal3 s 79200 70184 80800 70304 6 m_wbs_dat_o_10[16]
port 307 nsew signal input
rlabel metal3 s 79200 70864 80800 70984 6 m_wbs_dat_o_10[17]
port 308 nsew signal input
rlabel metal3 s 79200 71408 80800 71528 6 m_wbs_dat_o_10[18]
port 309 nsew signal input
rlabel metal3 s 79200 72088 80800 72208 6 m_wbs_dat_o_10[19]
port 310 nsew signal input
rlabel metal3 s 79200 60800 80800 60920 6 m_wbs_dat_o_10[1]
port 311 nsew signal input
rlabel metal3 s 79200 72632 80800 72752 6 m_wbs_dat_o_10[20]
port 312 nsew signal input
rlabel metal3 s 79200 73312 80800 73432 6 m_wbs_dat_o_10[21]
port 313 nsew signal input
rlabel metal3 s 79200 73992 80800 74112 6 m_wbs_dat_o_10[22]
port 314 nsew signal input
rlabel metal3 s 79200 74536 80800 74656 6 m_wbs_dat_o_10[23]
port 315 nsew signal input
rlabel metal3 s 79200 75216 80800 75336 6 m_wbs_dat_o_10[24]
port 316 nsew signal input
rlabel metal3 s 79200 75760 80800 75880 6 m_wbs_dat_o_10[25]
port 317 nsew signal input
rlabel metal3 s 79200 76440 80800 76560 6 m_wbs_dat_o_10[26]
port 318 nsew signal input
rlabel metal3 s 79200 77120 80800 77240 6 m_wbs_dat_o_10[27]
port 319 nsew signal input
rlabel metal3 s 79200 77664 80800 77784 6 m_wbs_dat_o_10[28]
port 320 nsew signal input
rlabel metal3 s 79200 78344 80800 78464 6 m_wbs_dat_o_10[29]
port 321 nsew signal input
rlabel metal3 s 79200 61480 80800 61600 6 m_wbs_dat_o_10[2]
port 322 nsew signal input
rlabel metal3 s 79200 78888 80800 79008 6 m_wbs_dat_o_10[30]
port 323 nsew signal input
rlabel metal3 s 79200 79568 80800 79688 6 m_wbs_dat_o_10[31]
port 324 nsew signal input
rlabel metal3 s 79200 62024 80800 62144 6 m_wbs_dat_o_10[3]
port 325 nsew signal input
rlabel metal3 s 79200 62704 80800 62824 6 m_wbs_dat_o_10[4]
port 326 nsew signal input
rlabel metal3 s 79200 63248 80800 63368 6 m_wbs_dat_o_10[5]
port 327 nsew signal input
rlabel metal3 s 79200 63928 80800 64048 6 m_wbs_dat_o_10[6]
port 328 nsew signal input
rlabel metal3 s 79200 64608 80800 64728 6 m_wbs_dat_o_10[7]
port 329 nsew signal input
rlabel metal3 s 79200 65152 80800 65272 6 m_wbs_dat_o_10[8]
port 330 nsew signal input
rlabel metal3 s 79200 65832 80800 65952 6 m_wbs_dat_o_10[9]
port 331 nsew signal input
rlabel metal3 s -800 41488 800 41608 4 m_wbs_dat_o_1[0]
port 332 nsew signal input
rlabel metal3 s -800 45432 800 45552 4 m_wbs_dat_o_1[10]
port 333 nsew signal input
rlabel metal3 s -800 45840 800 45960 4 m_wbs_dat_o_1[11]
port 334 nsew signal input
rlabel metal3 s -800 46248 800 46368 4 m_wbs_dat_o_1[12]
port 335 nsew signal input
rlabel metal3 s -800 46656 800 46776 4 m_wbs_dat_o_1[13]
port 336 nsew signal input
rlabel metal3 s -800 47064 800 47184 4 m_wbs_dat_o_1[14]
port 337 nsew signal input
rlabel metal3 s -800 47472 800 47592 4 m_wbs_dat_o_1[15]
port 338 nsew signal input
rlabel metal3 s -800 47880 800 48000 4 m_wbs_dat_o_1[16]
port 339 nsew signal input
rlabel metal3 s -800 48288 800 48408 4 m_wbs_dat_o_1[17]
port 340 nsew signal input
rlabel metal3 s -800 48696 800 48816 4 m_wbs_dat_o_1[18]
port 341 nsew signal input
rlabel metal3 s -800 49104 800 49224 4 m_wbs_dat_o_1[19]
port 342 nsew signal input
rlabel metal3 s -800 41896 800 42016 4 m_wbs_dat_o_1[1]
port 343 nsew signal input
rlabel metal3 s -800 49512 800 49632 4 m_wbs_dat_o_1[20]
port 344 nsew signal input
rlabel metal3 s -800 49920 800 50040 4 m_wbs_dat_o_1[21]
port 345 nsew signal input
rlabel metal3 s -800 50328 800 50448 4 m_wbs_dat_o_1[22]
port 346 nsew signal input
rlabel metal3 s -800 50736 800 50856 4 m_wbs_dat_o_1[23]
port 347 nsew signal input
rlabel metal3 s -800 51144 800 51264 4 m_wbs_dat_o_1[24]
port 348 nsew signal input
rlabel metal3 s -800 51552 800 51672 4 m_wbs_dat_o_1[25]
port 349 nsew signal input
rlabel metal3 s -800 51960 800 52080 4 m_wbs_dat_o_1[26]
port 350 nsew signal input
rlabel metal3 s -800 52368 800 52488 4 m_wbs_dat_o_1[27]
port 351 nsew signal input
rlabel metal3 s -800 52776 800 52896 4 m_wbs_dat_o_1[28]
port 352 nsew signal input
rlabel metal3 s -800 53184 800 53304 4 m_wbs_dat_o_1[29]
port 353 nsew signal input
rlabel metal3 s -800 42304 800 42424 4 m_wbs_dat_o_1[2]
port 354 nsew signal input
rlabel metal3 s -800 53456 800 53576 4 m_wbs_dat_o_1[30]
port 355 nsew signal input
rlabel metal3 s -800 53864 800 53984 4 m_wbs_dat_o_1[31]
port 356 nsew signal input
rlabel metal3 s -800 42712 800 42832 4 m_wbs_dat_o_1[3]
port 357 nsew signal input
rlabel metal3 s -800 43120 800 43240 4 m_wbs_dat_o_1[4]
port 358 nsew signal input
rlabel metal3 s -800 43528 800 43648 4 m_wbs_dat_o_1[5]
port 359 nsew signal input
rlabel metal3 s -800 43936 800 44056 4 m_wbs_dat_o_1[6]
port 360 nsew signal input
rlabel metal3 s -800 44344 800 44464 4 m_wbs_dat_o_1[7]
port 361 nsew signal input
rlabel metal3 s -800 44616 800 44736 4 m_wbs_dat_o_1[8]
port 362 nsew signal input
rlabel metal3 s -800 45024 800 45144 4 m_wbs_dat_o_1[9]
port 363 nsew signal input
rlabel metal3 s -800 54272 800 54392 4 m_wbs_dat_o_2[0]
port 364 nsew signal input
rlabel metal3 s -800 58352 800 58472 4 m_wbs_dat_o_2[10]
port 365 nsew signal input
rlabel metal3 s -800 58760 800 58880 4 m_wbs_dat_o_2[11]
port 366 nsew signal input
rlabel metal3 s -800 59168 800 59288 4 m_wbs_dat_o_2[12]
port 367 nsew signal input
rlabel metal3 s -800 59576 800 59696 4 m_wbs_dat_o_2[13]
port 368 nsew signal input
rlabel metal3 s -800 59984 800 60104 4 m_wbs_dat_o_2[14]
port 369 nsew signal input
rlabel metal3 s -800 60392 800 60512 4 m_wbs_dat_o_2[15]
port 370 nsew signal input
rlabel metal3 s -800 60800 800 60920 4 m_wbs_dat_o_2[16]
port 371 nsew signal input
rlabel metal3 s -800 61208 800 61328 4 m_wbs_dat_o_2[17]
port 372 nsew signal input
rlabel metal3 s -800 61616 800 61736 4 m_wbs_dat_o_2[18]
port 373 nsew signal input
rlabel metal3 s -800 62024 800 62144 4 m_wbs_dat_o_2[19]
port 374 nsew signal input
rlabel metal3 s -800 54680 800 54800 4 m_wbs_dat_o_2[1]
port 375 nsew signal input
rlabel metal3 s -800 62296 800 62416 4 m_wbs_dat_o_2[20]
port 376 nsew signal input
rlabel metal3 s -800 62704 800 62824 4 m_wbs_dat_o_2[21]
port 377 nsew signal input
rlabel metal3 s -800 63112 800 63232 4 m_wbs_dat_o_2[22]
port 378 nsew signal input
rlabel metal3 s -800 63520 800 63640 4 m_wbs_dat_o_2[23]
port 379 nsew signal input
rlabel metal3 s -800 63928 800 64048 4 m_wbs_dat_o_2[24]
port 380 nsew signal input
rlabel metal3 s -800 64336 800 64456 4 m_wbs_dat_o_2[25]
port 381 nsew signal input
rlabel metal3 s -800 64744 800 64864 4 m_wbs_dat_o_2[26]
port 382 nsew signal input
rlabel metal3 s -800 65152 800 65272 4 m_wbs_dat_o_2[27]
port 383 nsew signal input
rlabel metal3 s -800 65560 800 65680 4 m_wbs_dat_o_2[28]
port 384 nsew signal input
rlabel metal3 s -800 65968 800 66088 4 m_wbs_dat_o_2[29]
port 385 nsew signal input
rlabel metal3 s -800 55088 800 55208 4 m_wbs_dat_o_2[2]
port 386 nsew signal input
rlabel metal3 s -800 66376 800 66496 4 m_wbs_dat_o_2[30]
port 387 nsew signal input
rlabel metal3 s -800 66784 800 66904 4 m_wbs_dat_o_2[31]
port 388 nsew signal input
rlabel metal3 s -800 55496 800 55616 4 m_wbs_dat_o_2[3]
port 389 nsew signal input
rlabel metal3 s -800 55904 800 56024 4 m_wbs_dat_o_2[4]
port 390 nsew signal input
rlabel metal3 s -800 56312 800 56432 4 m_wbs_dat_o_2[5]
port 391 nsew signal input
rlabel metal3 s -800 56720 800 56840 4 m_wbs_dat_o_2[6]
port 392 nsew signal input
rlabel metal3 s -800 57128 800 57248 4 m_wbs_dat_o_2[7]
port 393 nsew signal input
rlabel metal3 s -800 57536 800 57656 4 m_wbs_dat_o_2[8]
port 394 nsew signal input
rlabel metal3 s -800 57944 800 58064 4 m_wbs_dat_o_2[9]
port 395 nsew signal input
rlabel metal3 s -800 67192 800 67312 4 m_wbs_dat_o_3[0]
port 396 nsew signal input
rlabel metal3 s -800 71136 800 71256 4 m_wbs_dat_o_3[10]
port 397 nsew signal input
rlabel metal3 s -800 71544 800 71664 4 m_wbs_dat_o_3[11]
port 398 nsew signal input
rlabel metal3 s -800 71952 800 72072 4 m_wbs_dat_o_3[12]
port 399 nsew signal input
rlabel metal3 s -800 72360 800 72480 4 m_wbs_dat_o_3[13]
port 400 nsew signal input
rlabel metal3 s -800 72768 800 72888 4 m_wbs_dat_o_3[14]
port 401 nsew signal input
rlabel metal3 s -800 73176 800 73296 4 m_wbs_dat_o_3[15]
port 402 nsew signal input
rlabel metal3 s -800 73584 800 73704 4 m_wbs_dat_o_3[16]
port 403 nsew signal input
rlabel metal3 s -800 73992 800 74112 4 m_wbs_dat_o_3[17]
port 404 nsew signal input
rlabel metal3 s -800 74400 800 74520 4 m_wbs_dat_o_3[18]
port 405 nsew signal input
rlabel metal3 s -800 74808 800 74928 4 m_wbs_dat_o_3[19]
port 406 nsew signal input
rlabel metal3 s -800 67600 800 67720 4 m_wbs_dat_o_3[1]
port 407 nsew signal input
rlabel metal3 s -800 75216 800 75336 4 m_wbs_dat_o_3[20]
port 408 nsew signal input
rlabel metal3 s -800 75624 800 75744 4 m_wbs_dat_o_3[21]
port 409 nsew signal input
rlabel metal3 s -800 76032 800 76152 4 m_wbs_dat_o_3[22]
port 410 nsew signal input
rlabel metal3 s -800 76440 800 76560 4 m_wbs_dat_o_3[23]
port 411 nsew signal input
rlabel metal3 s -800 76848 800 76968 4 m_wbs_dat_o_3[24]
port 412 nsew signal input
rlabel metal3 s -800 77256 800 77376 4 m_wbs_dat_o_3[25]
port 413 nsew signal input
rlabel metal3 s -800 77664 800 77784 4 m_wbs_dat_o_3[26]
port 414 nsew signal input
rlabel metal3 s -800 78072 800 78192 4 m_wbs_dat_o_3[27]
port 415 nsew signal input
rlabel metal3 s -800 78480 800 78600 4 m_wbs_dat_o_3[28]
port 416 nsew signal input
rlabel metal3 s -800 78888 800 79008 4 m_wbs_dat_o_3[29]
port 417 nsew signal input
rlabel metal3 s -800 68008 800 68128 4 m_wbs_dat_o_3[2]
port 418 nsew signal input
rlabel metal3 s -800 79296 800 79416 4 m_wbs_dat_o_3[30]
port 419 nsew signal input
rlabel metal3 s -800 79704 800 79824 4 m_wbs_dat_o_3[31]
port 420 nsew signal input
rlabel metal3 s -800 68416 800 68536 4 m_wbs_dat_o_3[3]
port 421 nsew signal input
rlabel metal3 s -800 68824 800 68944 4 m_wbs_dat_o_3[4]
port 422 nsew signal input
rlabel metal3 s -800 69232 800 69352 4 m_wbs_dat_o_3[5]
port 423 nsew signal input
rlabel metal3 s -800 69640 800 69760 4 m_wbs_dat_o_3[6]
port 424 nsew signal input
rlabel metal3 s -800 70048 800 70168 4 m_wbs_dat_o_3[7]
port 425 nsew signal input
rlabel metal3 s -800 70456 800 70576 4 m_wbs_dat_o_3[8]
port 426 nsew signal input
rlabel metal3 s -800 70864 800 70984 4 m_wbs_dat_o_3[9]
port 427 nsew signal input
rlabel metal2 s 48502 79200 48558 80800 6 m_wbs_dat_o_4[0]
port 428 nsew signal input
rlabel metal2 s 51814 79200 51870 80800 6 m_wbs_dat_o_4[10]
port 429 nsew signal input
rlabel metal2 s 52090 79200 52146 80800 6 m_wbs_dat_o_4[11]
port 430 nsew signal input
rlabel metal2 s 52458 79200 52514 80800 6 m_wbs_dat_o_4[12]
port 431 nsew signal input
rlabel metal2 s 52734 79200 52790 80800 6 m_wbs_dat_o_4[13]
port 432 nsew signal input
rlabel metal2 s 53102 79200 53158 80800 6 m_wbs_dat_o_4[14]
port 433 nsew signal input
rlabel metal2 s 53470 79200 53526 80800 6 m_wbs_dat_o_4[15]
port 434 nsew signal input
rlabel metal2 s 53746 79200 53802 80800 6 m_wbs_dat_o_4[16]
port 435 nsew signal input
rlabel metal2 s 54114 79200 54170 80800 6 m_wbs_dat_o_4[17]
port 436 nsew signal input
rlabel metal2 s 54390 79200 54446 80800 6 m_wbs_dat_o_4[18]
port 437 nsew signal input
rlabel metal2 s 54758 79200 54814 80800 6 m_wbs_dat_o_4[19]
port 438 nsew signal input
rlabel metal2 s 48778 79200 48834 80800 6 m_wbs_dat_o_4[1]
port 439 nsew signal input
rlabel metal2 s 55034 79200 55090 80800 6 m_wbs_dat_o_4[20]
port 440 nsew signal input
rlabel metal2 s 55402 79200 55458 80800 6 m_wbs_dat_o_4[21]
port 441 nsew signal input
rlabel metal2 s 55770 79200 55826 80800 6 m_wbs_dat_o_4[22]
port 442 nsew signal input
rlabel metal2 s 56046 79200 56102 80800 6 m_wbs_dat_o_4[23]
port 443 nsew signal input
rlabel metal2 s 56414 79200 56470 80800 6 m_wbs_dat_o_4[24]
port 444 nsew signal input
rlabel metal2 s 56690 79200 56746 80800 6 m_wbs_dat_o_4[25]
port 445 nsew signal input
rlabel metal2 s 57058 79200 57114 80800 6 m_wbs_dat_o_4[26]
port 446 nsew signal input
rlabel metal2 s 57334 79200 57390 80800 6 m_wbs_dat_o_4[27]
port 447 nsew signal input
rlabel metal2 s 57702 79200 57758 80800 6 m_wbs_dat_o_4[28]
port 448 nsew signal input
rlabel metal2 s 58070 79200 58126 80800 6 m_wbs_dat_o_4[29]
port 449 nsew signal input
rlabel metal2 s 49146 79200 49202 80800 6 m_wbs_dat_o_4[2]
port 450 nsew signal input
rlabel metal2 s 58346 79200 58402 80800 6 m_wbs_dat_o_4[30]
port 451 nsew signal input
rlabel metal2 s 58714 79200 58770 80800 6 m_wbs_dat_o_4[31]
port 452 nsew signal input
rlabel metal2 s 49514 79200 49570 80800 6 m_wbs_dat_o_4[3]
port 453 nsew signal input
rlabel metal2 s 49790 79200 49846 80800 6 m_wbs_dat_o_4[4]
port 454 nsew signal input
rlabel metal2 s 50158 79200 50214 80800 6 m_wbs_dat_o_4[5]
port 455 nsew signal input
rlabel metal2 s 50434 79200 50490 80800 6 m_wbs_dat_o_4[6]
port 456 nsew signal input
rlabel metal2 s 50802 79200 50858 80800 6 m_wbs_dat_o_4[7]
port 457 nsew signal input
rlabel metal2 s 51078 79200 51134 80800 6 m_wbs_dat_o_4[8]
port 458 nsew signal input
rlabel metal2 s 51446 79200 51502 80800 6 m_wbs_dat_o_4[9]
port 459 nsew signal input
rlabel metal2 s 58990 79200 59046 80800 6 m_wbs_dat_o_5[0]
port 460 nsew signal input
rlabel metal2 s 62302 79200 62358 80800 6 m_wbs_dat_o_5[10]
port 461 nsew signal input
rlabel metal2 s 62670 79200 62726 80800 6 m_wbs_dat_o_5[11]
port 462 nsew signal input
rlabel metal2 s 62946 79200 63002 80800 6 m_wbs_dat_o_5[12]
port 463 nsew signal input
rlabel metal2 s 63314 79200 63370 80800 6 m_wbs_dat_o_5[13]
port 464 nsew signal input
rlabel metal2 s 63590 79200 63646 80800 6 m_wbs_dat_o_5[14]
port 465 nsew signal input
rlabel metal2 s 63958 79200 64014 80800 6 m_wbs_dat_o_5[15]
port 466 nsew signal input
rlabel metal2 s 64326 79200 64382 80800 6 m_wbs_dat_o_5[16]
port 467 nsew signal input
rlabel metal2 s 64602 79200 64658 80800 6 m_wbs_dat_o_5[17]
port 468 nsew signal input
rlabel metal2 s 64970 79200 65026 80800 6 m_wbs_dat_o_5[18]
port 469 nsew signal input
rlabel metal2 s 65246 79200 65302 80800 6 m_wbs_dat_o_5[19]
port 470 nsew signal input
rlabel metal2 s 59358 79200 59414 80800 6 m_wbs_dat_o_5[1]
port 471 nsew signal input
rlabel metal2 s 65614 79200 65670 80800 6 m_wbs_dat_o_5[20]
port 472 nsew signal input
rlabel metal2 s 65982 79200 66038 80800 6 m_wbs_dat_o_5[21]
port 473 nsew signal input
rlabel metal2 s 66258 79200 66314 80800 6 m_wbs_dat_o_5[22]
port 474 nsew signal input
rlabel metal2 s 66626 79200 66682 80800 6 m_wbs_dat_o_5[23]
port 475 nsew signal input
rlabel metal2 s 66902 79200 66958 80800 6 m_wbs_dat_o_5[24]
port 476 nsew signal input
rlabel metal2 s 67270 79200 67326 80800 6 m_wbs_dat_o_5[25]
port 477 nsew signal input
rlabel metal2 s 67546 79200 67602 80800 6 m_wbs_dat_o_5[26]
port 478 nsew signal input
rlabel metal2 s 67914 79200 67970 80800 6 m_wbs_dat_o_5[27]
port 479 nsew signal input
rlabel metal2 s 68282 79200 68338 80800 6 m_wbs_dat_o_5[28]
port 480 nsew signal input
rlabel metal2 s 68558 79200 68614 80800 6 m_wbs_dat_o_5[29]
port 481 nsew signal input
rlabel metal2 s 59726 79200 59782 80800 6 m_wbs_dat_o_5[2]
port 482 nsew signal input
rlabel metal2 s 68926 79200 68982 80800 6 m_wbs_dat_o_5[30]
port 483 nsew signal input
rlabel metal2 s 69202 79200 69258 80800 6 m_wbs_dat_o_5[31]
port 484 nsew signal input
rlabel metal2 s 60002 79200 60058 80800 6 m_wbs_dat_o_5[3]
port 485 nsew signal input
rlabel metal2 s 60370 79200 60426 80800 6 m_wbs_dat_o_5[4]
port 486 nsew signal input
rlabel metal2 s 60646 79200 60702 80800 6 m_wbs_dat_o_5[5]
port 487 nsew signal input
rlabel metal2 s 61014 79200 61070 80800 6 m_wbs_dat_o_5[6]
port 488 nsew signal input
rlabel metal2 s 61290 79200 61346 80800 6 m_wbs_dat_o_5[7]
port 489 nsew signal input
rlabel metal2 s 61658 79200 61714 80800 6 m_wbs_dat_o_5[8]
port 490 nsew signal input
rlabel metal2 s 62026 79200 62082 80800 6 m_wbs_dat_o_5[9]
port 491 nsew signal input
rlabel metal2 s 69570 79200 69626 80800 6 m_wbs_dat_o_6[0]
port 492 nsew signal input
rlabel metal2 s 72882 79200 72938 80800 6 m_wbs_dat_o_6[10]
port 493 nsew signal input
rlabel metal2 s 73158 79200 73214 80800 6 m_wbs_dat_o_6[11]
port 494 nsew signal input
rlabel metal2 s 73526 79200 73582 80800 6 m_wbs_dat_o_6[12]
port 495 nsew signal input
rlabel metal2 s 73802 79200 73858 80800 6 m_wbs_dat_o_6[13]
port 496 nsew signal input
rlabel metal2 s 74170 79200 74226 80800 6 m_wbs_dat_o_6[14]
port 497 nsew signal input
rlabel metal2 s 74538 79200 74594 80800 6 m_wbs_dat_o_6[15]
port 498 nsew signal input
rlabel metal2 s 74814 79200 74870 80800 6 m_wbs_dat_o_6[16]
port 499 nsew signal input
rlabel metal2 s 75182 79200 75238 80800 6 m_wbs_dat_o_6[17]
port 500 nsew signal input
rlabel metal2 s 75458 79200 75514 80800 6 m_wbs_dat_o_6[18]
port 501 nsew signal input
rlabel metal2 s 75826 79200 75882 80800 6 m_wbs_dat_o_6[19]
port 502 nsew signal input
rlabel metal2 s 69938 79200 69994 80800 6 m_wbs_dat_o_6[1]
port 503 nsew signal input
rlabel metal2 s 76194 79200 76250 80800 6 m_wbs_dat_o_6[20]
port 504 nsew signal input
rlabel metal2 s 76470 79200 76526 80800 6 m_wbs_dat_o_6[21]
port 505 nsew signal input
rlabel metal2 s 76838 79200 76894 80800 6 m_wbs_dat_o_6[22]
port 506 nsew signal input
rlabel metal2 s 77114 79200 77170 80800 6 m_wbs_dat_o_6[23]
port 507 nsew signal input
rlabel metal2 s 77482 79200 77538 80800 6 m_wbs_dat_o_6[24]
port 508 nsew signal input
rlabel metal2 s 77758 79200 77814 80800 6 m_wbs_dat_o_6[25]
port 509 nsew signal input
rlabel metal2 s 78126 79200 78182 80800 6 m_wbs_dat_o_6[26]
port 510 nsew signal input
rlabel metal2 s 78494 79200 78550 80800 6 m_wbs_dat_o_6[27]
port 511 nsew signal input
rlabel metal2 s 78770 79200 78826 80800 6 m_wbs_dat_o_6[28]
port 512 nsew signal input
rlabel metal2 s 79138 79200 79194 80800 6 m_wbs_dat_o_6[29]
port 513 nsew signal input
rlabel metal2 s 70214 79200 70270 80800 6 m_wbs_dat_o_6[2]
port 514 nsew signal input
rlabel metal2 s 79414 79200 79470 80800 6 m_wbs_dat_o_6[30]
port 515 nsew signal input
rlabel metal2 s 79782 79200 79838 80800 6 m_wbs_dat_o_6[31]
port 516 nsew signal input
rlabel metal2 s 70582 79200 70638 80800 6 m_wbs_dat_o_6[3]
port 517 nsew signal input
rlabel metal2 s 70858 79200 70914 80800 6 m_wbs_dat_o_6[4]
port 518 nsew signal input
rlabel metal2 s 71226 79200 71282 80800 6 m_wbs_dat_o_6[5]
port 519 nsew signal input
rlabel metal2 s 71502 79200 71558 80800 6 m_wbs_dat_o_6[6]
port 520 nsew signal input
rlabel metal2 s 71870 79200 71926 80800 6 m_wbs_dat_o_6[7]
port 521 nsew signal input
rlabel metal2 s 72238 79200 72294 80800 6 m_wbs_dat_o_6[8]
port 522 nsew signal input
rlabel metal2 s 72514 79200 72570 80800 6 m_wbs_dat_o_6[9]
port 523 nsew signal input
rlabel metal3 s 79200 280 80800 400 6 m_wbs_dat_o_7[0]
port 524 nsew signal input
rlabel metal3 s 79200 6400 80800 6520 6 m_wbs_dat_o_7[10]
port 525 nsew signal input
rlabel metal3 s 79200 7080 80800 7200 6 m_wbs_dat_o_7[11]
port 526 nsew signal input
rlabel metal3 s 79200 7760 80800 7880 6 m_wbs_dat_o_7[12]
port 527 nsew signal input
rlabel metal3 s 79200 8304 80800 8424 6 m_wbs_dat_o_7[13]
port 528 nsew signal input
rlabel metal3 s 79200 8984 80800 9104 6 m_wbs_dat_o_7[14]
port 529 nsew signal input
rlabel metal3 s 79200 9528 80800 9648 6 m_wbs_dat_o_7[15]
port 530 nsew signal input
rlabel metal3 s 79200 10208 80800 10328 6 m_wbs_dat_o_7[16]
port 531 nsew signal input
rlabel metal3 s 79200 10888 80800 11008 6 m_wbs_dat_o_7[17]
port 532 nsew signal input
rlabel metal3 s 79200 11432 80800 11552 6 m_wbs_dat_o_7[18]
port 533 nsew signal input
rlabel metal3 s 79200 12112 80800 12232 6 m_wbs_dat_o_7[19]
port 534 nsew signal input
rlabel metal3 s 79200 824 80800 944 6 m_wbs_dat_o_7[1]
port 535 nsew signal input
rlabel metal3 s 79200 12656 80800 12776 6 m_wbs_dat_o_7[20]
port 536 nsew signal input
rlabel metal3 s 79200 13336 80800 13456 6 m_wbs_dat_o_7[21]
port 537 nsew signal input
rlabel metal3 s 79200 14016 80800 14136 6 m_wbs_dat_o_7[22]
port 538 nsew signal input
rlabel metal3 s 79200 14560 80800 14680 6 m_wbs_dat_o_7[23]
port 539 nsew signal input
rlabel metal3 s 79200 15240 80800 15360 6 m_wbs_dat_o_7[24]
port 540 nsew signal input
rlabel metal3 s 79200 15784 80800 15904 6 m_wbs_dat_o_7[25]
port 541 nsew signal input
rlabel metal3 s 79200 16464 80800 16584 6 m_wbs_dat_o_7[26]
port 542 nsew signal input
rlabel metal3 s 79200 17144 80800 17264 6 m_wbs_dat_o_7[27]
port 543 nsew signal input
rlabel metal3 s 79200 17688 80800 17808 6 m_wbs_dat_o_7[28]
port 544 nsew signal input
rlabel metal3 s 79200 18368 80800 18488 6 m_wbs_dat_o_7[29]
port 545 nsew signal input
rlabel metal3 s 79200 1504 80800 1624 6 m_wbs_dat_o_7[2]
port 546 nsew signal input
rlabel metal3 s 79200 18912 80800 19032 6 m_wbs_dat_o_7[30]
port 547 nsew signal input
rlabel metal3 s 79200 19592 80800 19712 6 m_wbs_dat_o_7[31]
port 548 nsew signal input
rlabel metal3 s 79200 2048 80800 2168 6 m_wbs_dat_o_7[3]
port 549 nsew signal input
rlabel metal3 s 79200 2728 80800 2848 6 m_wbs_dat_o_7[4]
port 550 nsew signal input
rlabel metal3 s 79200 3272 80800 3392 6 m_wbs_dat_o_7[5]
port 551 nsew signal input
rlabel metal3 s 79200 3952 80800 4072 6 m_wbs_dat_o_7[6]
port 552 nsew signal input
rlabel metal3 s 79200 4632 80800 4752 6 m_wbs_dat_o_7[7]
port 553 nsew signal input
rlabel metal3 s 79200 5176 80800 5296 6 m_wbs_dat_o_7[8]
port 554 nsew signal input
rlabel metal3 s 79200 5856 80800 5976 6 m_wbs_dat_o_7[9]
port 555 nsew signal input
rlabel metal3 s 79200 20272 80800 20392 6 m_wbs_dat_o_8[0]
port 556 nsew signal input
rlabel metal3 s 79200 26392 80800 26512 6 m_wbs_dat_o_8[10]
port 557 nsew signal input
rlabel metal3 s 79200 27072 80800 27192 6 m_wbs_dat_o_8[11]
port 558 nsew signal input
rlabel metal3 s 79200 27752 80800 27872 6 m_wbs_dat_o_8[12]
port 559 nsew signal input
rlabel metal3 s 79200 28296 80800 28416 6 m_wbs_dat_o_8[13]
port 560 nsew signal input
rlabel metal3 s 79200 28976 80800 29096 6 m_wbs_dat_o_8[14]
port 561 nsew signal input
rlabel metal3 s 79200 29520 80800 29640 6 m_wbs_dat_o_8[15]
port 562 nsew signal input
rlabel metal3 s 79200 30200 80800 30320 6 m_wbs_dat_o_8[16]
port 563 nsew signal input
rlabel metal3 s 79200 30880 80800 31000 6 m_wbs_dat_o_8[17]
port 564 nsew signal input
rlabel metal3 s 79200 31424 80800 31544 6 m_wbs_dat_o_8[18]
port 565 nsew signal input
rlabel metal3 s 79200 32104 80800 32224 6 m_wbs_dat_o_8[19]
port 566 nsew signal input
rlabel metal3 s 79200 20816 80800 20936 6 m_wbs_dat_o_8[1]
port 567 nsew signal input
rlabel metal3 s 79200 32648 80800 32768 6 m_wbs_dat_o_8[20]
port 568 nsew signal input
rlabel metal3 s 79200 33328 80800 33448 6 m_wbs_dat_o_8[21]
port 569 nsew signal input
rlabel metal3 s 79200 34008 80800 34128 6 m_wbs_dat_o_8[22]
port 570 nsew signal input
rlabel metal3 s 79200 34552 80800 34672 6 m_wbs_dat_o_8[23]
port 571 nsew signal input
rlabel metal3 s 79200 35232 80800 35352 6 m_wbs_dat_o_8[24]
port 572 nsew signal input
rlabel metal3 s 79200 35776 80800 35896 6 m_wbs_dat_o_8[25]
port 573 nsew signal input
rlabel metal3 s 79200 36456 80800 36576 6 m_wbs_dat_o_8[26]
port 574 nsew signal input
rlabel metal3 s 79200 37136 80800 37256 6 m_wbs_dat_o_8[27]
port 575 nsew signal input
rlabel metal3 s 79200 37680 80800 37800 6 m_wbs_dat_o_8[28]
port 576 nsew signal input
rlabel metal3 s 79200 38360 80800 38480 6 m_wbs_dat_o_8[29]
port 577 nsew signal input
rlabel metal3 s 79200 21496 80800 21616 6 m_wbs_dat_o_8[2]
port 578 nsew signal input
rlabel metal3 s 79200 38904 80800 39024 6 m_wbs_dat_o_8[30]
port 579 nsew signal input
rlabel metal3 s 79200 39584 80800 39704 6 m_wbs_dat_o_8[31]
port 580 nsew signal input
rlabel metal3 s 79200 22040 80800 22160 6 m_wbs_dat_o_8[3]
port 581 nsew signal input
rlabel metal3 s 79200 22720 80800 22840 6 m_wbs_dat_o_8[4]
port 582 nsew signal input
rlabel metal3 s 79200 23264 80800 23384 6 m_wbs_dat_o_8[5]
port 583 nsew signal input
rlabel metal3 s 79200 23944 80800 24064 6 m_wbs_dat_o_8[6]
port 584 nsew signal input
rlabel metal3 s 79200 24624 80800 24744 6 m_wbs_dat_o_8[7]
port 585 nsew signal input
rlabel metal3 s 79200 25168 80800 25288 6 m_wbs_dat_o_8[8]
port 586 nsew signal input
rlabel metal3 s 79200 25848 80800 25968 6 m_wbs_dat_o_8[9]
port 587 nsew signal input
rlabel metal3 s 79200 40264 80800 40384 6 m_wbs_dat_o_9[0]
port 588 nsew signal input
rlabel metal3 s 79200 46384 80800 46504 6 m_wbs_dat_o_9[10]
port 589 nsew signal input
rlabel metal3 s 79200 47064 80800 47184 6 m_wbs_dat_o_9[11]
port 590 nsew signal input
rlabel metal3 s 79200 47744 80800 47864 6 m_wbs_dat_o_9[12]
port 591 nsew signal input
rlabel metal3 s 79200 48288 80800 48408 6 m_wbs_dat_o_9[13]
port 592 nsew signal input
rlabel metal3 s 79200 48968 80800 49088 6 m_wbs_dat_o_9[14]
port 593 nsew signal input
rlabel metal3 s 79200 49512 80800 49632 6 m_wbs_dat_o_9[15]
port 594 nsew signal input
rlabel metal3 s 79200 50192 80800 50312 6 m_wbs_dat_o_9[16]
port 595 nsew signal input
rlabel metal3 s 79200 50872 80800 50992 6 m_wbs_dat_o_9[17]
port 596 nsew signal input
rlabel metal3 s 79200 51416 80800 51536 6 m_wbs_dat_o_9[18]
port 597 nsew signal input
rlabel metal3 s 79200 52096 80800 52216 6 m_wbs_dat_o_9[19]
port 598 nsew signal input
rlabel metal3 s 79200 40808 80800 40928 6 m_wbs_dat_o_9[1]
port 599 nsew signal input
rlabel metal3 s 79200 52640 80800 52760 6 m_wbs_dat_o_9[20]
port 600 nsew signal input
rlabel metal3 s 79200 53320 80800 53440 6 m_wbs_dat_o_9[21]
port 601 nsew signal input
rlabel metal3 s 79200 54000 80800 54120 6 m_wbs_dat_o_9[22]
port 602 nsew signal input
rlabel metal3 s 79200 54544 80800 54664 6 m_wbs_dat_o_9[23]
port 603 nsew signal input
rlabel metal3 s 79200 55224 80800 55344 6 m_wbs_dat_o_9[24]
port 604 nsew signal input
rlabel metal3 s 79200 55768 80800 55888 6 m_wbs_dat_o_9[25]
port 605 nsew signal input
rlabel metal3 s 79200 56448 80800 56568 6 m_wbs_dat_o_9[26]
port 606 nsew signal input
rlabel metal3 s 79200 57128 80800 57248 6 m_wbs_dat_o_9[27]
port 607 nsew signal input
rlabel metal3 s 79200 57672 80800 57792 6 m_wbs_dat_o_9[28]
port 608 nsew signal input
rlabel metal3 s 79200 58352 80800 58472 6 m_wbs_dat_o_9[29]
port 609 nsew signal input
rlabel metal3 s 79200 41488 80800 41608 6 m_wbs_dat_o_9[2]
port 610 nsew signal input
rlabel metal3 s 79200 58896 80800 59016 6 m_wbs_dat_o_9[30]
port 611 nsew signal input
rlabel metal3 s 79200 59576 80800 59696 6 m_wbs_dat_o_9[31]
port 612 nsew signal input
rlabel metal3 s 79200 42032 80800 42152 6 m_wbs_dat_o_9[3]
port 613 nsew signal input
rlabel metal3 s 79200 42712 80800 42832 6 m_wbs_dat_o_9[4]
port 614 nsew signal input
rlabel metal3 s 79200 43256 80800 43376 6 m_wbs_dat_o_9[5]
port 615 nsew signal input
rlabel metal3 s 79200 43936 80800 44056 6 m_wbs_dat_o_9[6]
port 616 nsew signal input
rlabel metal3 s 79200 44616 80800 44736 6 m_wbs_dat_o_9[7]
port 617 nsew signal input
rlabel metal3 s 79200 45160 80800 45280 6 m_wbs_dat_o_9[8]
port 618 nsew signal input
rlabel metal3 s 79200 45840 80800 45960 6 m_wbs_dat_o_9[9]
port 619 nsew signal input
rlabel metal2 s 41234 79200 41290 80800 6 m_wbs_stb_i[0]
port 620 nsew signal output
rlabel metal2 s 44546 79200 44602 80800 6 m_wbs_stb_i[10]
port 621 nsew signal output
rlabel metal2 s 41602 79200 41658 80800 6 m_wbs_stb_i[1]
port 622 nsew signal output
rlabel metal2 s 41878 79200 41934 80800 6 m_wbs_stb_i[2]
port 623 nsew signal output
rlabel metal2 s 42246 79200 42302 80800 6 m_wbs_stb_i[3]
port 624 nsew signal output
rlabel metal2 s 42522 79200 42578 80800 6 m_wbs_stb_i[4]
port 625 nsew signal output
rlabel metal2 s 42890 79200 42946 80800 6 m_wbs_stb_i[5]
port 626 nsew signal output
rlabel metal2 s 43258 79200 43314 80800 6 m_wbs_stb_i[6]
port 627 nsew signal output
rlabel metal2 s 43534 79200 43590 80800 6 m_wbs_stb_i[7]
port 628 nsew signal output
rlabel metal2 s 43902 79200 43958 80800 6 m_wbs_stb_i[8]
port 629 nsew signal output
rlabel metal2 s 44178 79200 44234 80800 6 m_wbs_stb_i[9]
port 630 nsew signal output
rlabel metal3 s -800 144 800 264 4 wb_clk_i
port 631 nsew signal input
rlabel metal3 s -800 416 800 536 4 wb_rst_i
port 632 nsew signal input
rlabel metal3 s -800 14152 800 14272 4 wbs_ack_o
port 633 nsew signal output
rlabel metal3 s -800 1232 800 1352 4 wbs_adr_i[0]
port 634 nsew signal input
rlabel metal3 s -800 5312 800 5432 4 wbs_adr_i[10]
port 635 nsew signal input
rlabel metal3 s -800 5720 800 5840 4 wbs_adr_i[11]
port 636 nsew signal input
rlabel metal3 s -800 6128 800 6248 4 wbs_adr_i[12]
port 637 nsew signal input
rlabel metal3 s -800 6536 800 6656 4 wbs_adr_i[13]
port 638 nsew signal input
rlabel metal3 s -800 6944 800 7064 4 wbs_adr_i[14]
port 639 nsew signal input
rlabel metal3 s -800 7352 800 7472 4 wbs_adr_i[15]
port 640 nsew signal input
rlabel metal3 s -800 7760 800 7880 4 wbs_adr_i[16]
port 641 nsew signal input
rlabel metal3 s -800 8168 800 8288 4 wbs_adr_i[17]
port 642 nsew signal input
rlabel metal3 s -800 8576 800 8696 4 wbs_adr_i[18]
port 643 nsew signal input
rlabel metal3 s -800 8984 800 9104 4 wbs_adr_i[19]
port 644 nsew signal input
rlabel metal3 s -800 1640 800 1760 4 wbs_adr_i[1]
port 645 nsew signal input
rlabel metal3 s -800 9256 800 9376 4 wbs_adr_i[20]
port 646 nsew signal input
rlabel metal3 s -800 9664 800 9784 4 wbs_adr_i[21]
port 647 nsew signal input
rlabel metal3 s -800 10072 800 10192 4 wbs_adr_i[22]
port 648 nsew signal input
rlabel metal3 s -800 10480 800 10600 4 wbs_adr_i[23]
port 649 nsew signal input
rlabel metal3 s -800 10888 800 11008 4 wbs_adr_i[24]
port 650 nsew signal input
rlabel metal3 s -800 11296 800 11416 4 wbs_adr_i[25]
port 651 nsew signal input
rlabel metal3 s -800 11704 800 11824 4 wbs_adr_i[26]
port 652 nsew signal input
rlabel metal3 s -800 12112 800 12232 4 wbs_adr_i[27]
port 653 nsew signal input
rlabel metal3 s -800 12520 800 12640 4 wbs_adr_i[28]
port 654 nsew signal input
rlabel metal3 s -800 12928 800 13048 4 wbs_adr_i[29]
port 655 nsew signal input
rlabel metal3 s -800 2048 800 2168 4 wbs_adr_i[2]
port 656 nsew signal input
rlabel metal3 s -800 13336 800 13456 4 wbs_adr_i[30]
port 657 nsew signal input
rlabel metal3 s -800 13744 800 13864 4 wbs_adr_i[31]
port 658 nsew signal input
rlabel metal3 s -800 2456 800 2576 4 wbs_adr_i[3]
port 659 nsew signal input
rlabel metal3 s -800 2864 800 2984 4 wbs_adr_i[4]
port 660 nsew signal input
rlabel metal3 s -800 3272 800 3392 4 wbs_adr_i[5]
port 661 nsew signal input
rlabel metal3 s -800 3680 800 3800 4 wbs_adr_i[6]
port 662 nsew signal input
rlabel metal3 s -800 4088 800 4208 4 wbs_adr_i[7]
port 663 nsew signal input
rlabel metal3 s -800 4496 800 4616 4 wbs_adr_i[8]
port 664 nsew signal input
rlabel metal3 s -800 4904 800 5024 4 wbs_adr_i[9]
port 665 nsew signal input
rlabel metal3 s -800 14560 800 14680 4 wbs_dat_o[0]
port 666 nsew signal output
rlabel metal3 s -800 18504 800 18624 4 wbs_dat_o[10]
port 667 nsew signal output
rlabel metal3 s -800 18912 800 19032 4 wbs_dat_o[11]
port 668 nsew signal output
rlabel metal3 s -800 19320 800 19440 4 wbs_dat_o[12]
port 669 nsew signal output
rlabel metal3 s -800 19728 800 19848 4 wbs_dat_o[13]
port 670 nsew signal output
rlabel metal3 s -800 20136 800 20256 4 wbs_dat_o[14]
port 671 nsew signal output
rlabel metal3 s -800 20544 800 20664 4 wbs_dat_o[15]
port 672 nsew signal output
rlabel metal3 s -800 20952 800 21072 4 wbs_dat_o[16]
port 673 nsew signal output
rlabel metal3 s -800 21360 800 21480 4 wbs_dat_o[17]
port 674 nsew signal output
rlabel metal3 s -800 21768 800 21888 4 wbs_dat_o[18]
port 675 nsew signal output
rlabel metal3 s -800 22176 800 22296 4 wbs_dat_o[19]
port 676 nsew signal output
rlabel metal3 s -800 14968 800 15088 4 wbs_dat_o[1]
port 677 nsew signal output
rlabel metal3 s -800 22584 800 22704 4 wbs_dat_o[20]
port 678 nsew signal output
rlabel metal3 s -800 22992 800 23112 4 wbs_dat_o[21]
port 679 nsew signal output
rlabel metal3 s -800 23400 800 23520 4 wbs_dat_o[22]
port 680 nsew signal output
rlabel metal3 s -800 23808 800 23928 4 wbs_dat_o[23]
port 681 nsew signal output
rlabel metal3 s -800 24216 800 24336 4 wbs_dat_o[24]
port 682 nsew signal output
rlabel metal3 s -800 24624 800 24744 4 wbs_dat_o[25]
port 683 nsew signal output
rlabel metal3 s -800 25032 800 25152 4 wbs_dat_o[26]
port 684 nsew signal output
rlabel metal3 s -800 25440 800 25560 4 wbs_dat_o[27]
port 685 nsew signal output
rlabel metal3 s -800 25848 800 25968 4 wbs_dat_o[28]
port 686 nsew signal output
rlabel metal3 s -800 26256 800 26376 4 wbs_dat_o[29]
port 687 nsew signal output
rlabel metal3 s -800 15376 800 15496 4 wbs_dat_o[2]
port 688 nsew signal output
rlabel metal3 s -800 26664 800 26784 4 wbs_dat_o[30]
port 689 nsew signal output
rlabel metal3 s -800 26936 800 27056 4 wbs_dat_o[31]
port 690 nsew signal output
rlabel metal3 s -800 15784 800 15904 4 wbs_dat_o[3]
port 691 nsew signal output
rlabel metal3 s -800 16192 800 16312 4 wbs_dat_o[4]
port 692 nsew signal output
rlabel metal3 s -800 16600 800 16720 4 wbs_dat_o[5]
port 693 nsew signal output
rlabel metal3 s -800 17008 800 17128 4 wbs_dat_o[6]
port 694 nsew signal output
rlabel metal3 s -800 17416 800 17536 4 wbs_dat_o[7]
port 695 nsew signal output
rlabel metal3 s -800 17824 800 17944 4 wbs_dat_o[8]
port 696 nsew signal output
rlabel metal3 s -800 18096 800 18216 4 wbs_dat_o[9]
port 697 nsew signal output
rlabel metal3 s -800 824 800 944 4 wbs_stb_i
port 698 nsew signal input
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 699 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 700 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 701 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 702 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 703 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 80000 80000
string LEFview TRUE
string GDS_FILE /project/openlane/multiplex/runs/multiplex/results/magic/multiplex.gds
string GDS_END 4893382
string GDS_START 219738
<< end >>

