module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    vccd2,
    vssd2,
    vdda1,
    vssa1,
    vdda2,
    vssa2,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 input vccd2;
 input vssd2;
 input vdda1;
 input vssa1;
 input vdda2;
 input vssa2;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 multiplex icon (.wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_stb_i(wbs_stb_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({io_in[37],
    io_in[36],
    io_in[35],
    io_in[34],
    io_in[33],
    io_in[32],
    io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21],
    io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .irq({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .la_data_in({la_data_in[10],
    la_data_in[9],
    la_data_in[8],
    la_data_in[7],
    la_data_in[6],
    la_data_in[5],
    la_data_in[4],
    la_data_in[3],
    la_data_in[2],
    la_data_in[1],
    la_data_in[0]}),
    .la_data_out({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96],
    la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64],
    la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .m_wb_rst_i({\m_wb_rst_i[10] ,
    \m_wb_rst_i[9] ,
    \m_wb_rst_i[8] ,
    \m_wb_rst_i[7] ,
    \m_wb_rst_i[6] ,
    \m_wb_rst_i[5] ,
    \m_wb_rst_i[4] ,
    \m_wb_rst_i[3] ,
    \m_wb_rst_i[2] ,
    \m_wb_rst_i[1] ,
    \m_wb_rst_i[0] }),
    .m_wbs_ack_o({\m_wbs_ack_out[10] ,
    \m_wbs_ack_out[9] ,
    \m_wbs_ack_out[8] ,
    \m_wbs_ack_out[7] ,
    \m_wbs_ack_out[6] ,
    \m_wbs_ack_out[5] ,
    \m_wbs_ack_out[4] ,
    \m_wbs_ack_out[3] ,
    \m_wbs_ack_out[2] ,
    \m_wbs_ack_out[1] ,
    \m_wbs_ack_out[0] }),
    .m_wbs_dat_o_0({\wbs_dat_out_0[31] ,
    \wbs_dat_out_0[30] ,
    \wbs_dat_out_0[29] ,
    \wbs_dat_out_0[28] ,
    \wbs_dat_out_0[27] ,
    \wbs_dat_out_0[26] ,
    \wbs_dat_out_0[25] ,
    \wbs_dat_out_0[24] ,
    \wbs_dat_out_0[23] ,
    \wbs_dat_out_0[22] ,
    \wbs_dat_out_0[21] ,
    \wbs_dat_out_0[20] ,
    \wbs_dat_out_0[19] ,
    \wbs_dat_out_0[18] ,
    \wbs_dat_out_0[17] ,
    \wbs_dat_out_0[16] ,
    \wbs_dat_out_0[15] ,
    \wbs_dat_out_0[14] ,
    \wbs_dat_out_0[13] ,
    \wbs_dat_out_0[12] ,
    \wbs_dat_out_0[11] ,
    \wbs_dat_out_0[10] ,
    \wbs_dat_out_0[9] ,
    \wbs_dat_out_0[8] ,
    \wbs_dat_out_0[7] ,
    \wbs_dat_out_0[6] ,
    \wbs_dat_out_0[5] ,
    \wbs_dat_out_0[4] ,
    \wbs_dat_out_0[3] ,
    \wbs_dat_out_0[2] ,
    \wbs_dat_out_0[1] ,
    \wbs_dat_out_0[0] }),
    .m_wbs_dat_o_1({\wbs_dat_out_1[31] ,
    \wbs_dat_out_1[30] ,
    \wbs_dat_out_1[29] ,
    \wbs_dat_out_1[28] ,
    \wbs_dat_out_1[27] ,
    \wbs_dat_out_1[26] ,
    \wbs_dat_out_1[25] ,
    \wbs_dat_out_1[24] ,
    \wbs_dat_out_1[23] ,
    \wbs_dat_out_1[22] ,
    \wbs_dat_out_1[21] ,
    \wbs_dat_out_1[20] ,
    \wbs_dat_out_1[19] ,
    \wbs_dat_out_1[18] ,
    \wbs_dat_out_1[17] ,
    \wbs_dat_out_1[16] ,
    \wbs_dat_out_1[15] ,
    \wbs_dat_out_1[14] ,
    \wbs_dat_out_1[13] ,
    \wbs_dat_out_1[12] ,
    \wbs_dat_out_1[11] ,
    \wbs_dat_out_1[10] ,
    \wbs_dat_out_1[9] ,
    \wbs_dat_out_1[8] ,
    \wbs_dat_out_1[7] ,
    \wbs_dat_out_1[6] ,
    \wbs_dat_out_1[5] ,
    \wbs_dat_out_1[4] ,
    \wbs_dat_out_1[3] ,
    \wbs_dat_out_1[2] ,
    \wbs_dat_out_1[1] ,
    \wbs_dat_out_1[0] }),
    .m_wbs_dat_o_10({\wbs_dat_out_10[31] ,
    \wbs_dat_out_10[30] ,
    \wbs_dat_out_10[29] ,
    \wbs_dat_out_10[28] ,
    \wbs_dat_out_10[27] ,
    \wbs_dat_out_10[26] ,
    \wbs_dat_out_10[25] ,
    \wbs_dat_out_10[24] ,
    \wbs_dat_out_10[23] ,
    \wbs_dat_out_10[22] ,
    \wbs_dat_out_10[21] ,
    \wbs_dat_out_10[20] ,
    \wbs_dat_out_10[19] ,
    \wbs_dat_out_10[18] ,
    \wbs_dat_out_10[17] ,
    \wbs_dat_out_10[16] ,
    \wbs_dat_out_10[15] ,
    \wbs_dat_out_10[14] ,
    \wbs_dat_out_10[13] ,
    \wbs_dat_out_10[12] ,
    \wbs_dat_out_10[11] ,
    \wbs_dat_out_10[10] ,
    \wbs_dat_out_10[9] ,
    \wbs_dat_out_10[8] ,
    \wbs_dat_out_10[7] ,
    \wbs_dat_out_10[6] ,
    \wbs_dat_out_10[5] ,
    \wbs_dat_out_10[4] ,
    \wbs_dat_out_10[3] ,
    \wbs_dat_out_10[2] ,
    \wbs_dat_out_10[1] ,
    \wbs_dat_out_10[0] }),
    .m_wbs_dat_o_2({\wbs_dat_out_2[31] ,
    \wbs_dat_out_2[30] ,
    \wbs_dat_out_2[29] ,
    \wbs_dat_out_2[28] ,
    \wbs_dat_out_2[27] ,
    \wbs_dat_out_2[26] ,
    \wbs_dat_out_2[25] ,
    \wbs_dat_out_2[24] ,
    \wbs_dat_out_2[23] ,
    \wbs_dat_out_2[22] ,
    \wbs_dat_out_2[21] ,
    \wbs_dat_out_2[20] ,
    \wbs_dat_out_2[19] ,
    \wbs_dat_out_2[18] ,
    \wbs_dat_out_2[17] ,
    \wbs_dat_out_2[16] ,
    \wbs_dat_out_2[15] ,
    \wbs_dat_out_2[14] ,
    \wbs_dat_out_2[13] ,
    \wbs_dat_out_2[12] ,
    \wbs_dat_out_2[11] ,
    \wbs_dat_out_2[10] ,
    \wbs_dat_out_2[9] ,
    \wbs_dat_out_2[8] ,
    \wbs_dat_out_2[7] ,
    \wbs_dat_out_2[6] ,
    \wbs_dat_out_2[5] ,
    \wbs_dat_out_2[4] ,
    \wbs_dat_out_2[3] ,
    \wbs_dat_out_2[2] ,
    \wbs_dat_out_2[1] ,
    \wbs_dat_out_2[0] }),
    .m_wbs_dat_o_3({\wbs_dat_out_3[31] ,
    \wbs_dat_out_3[30] ,
    \wbs_dat_out_3[29] ,
    \wbs_dat_out_3[28] ,
    \wbs_dat_out_3[27] ,
    \wbs_dat_out_3[26] ,
    \wbs_dat_out_3[25] ,
    \wbs_dat_out_3[24] ,
    \wbs_dat_out_3[23] ,
    \wbs_dat_out_3[22] ,
    \wbs_dat_out_3[21] ,
    \wbs_dat_out_3[20] ,
    \wbs_dat_out_3[19] ,
    \wbs_dat_out_3[18] ,
    \wbs_dat_out_3[17] ,
    \wbs_dat_out_3[16] ,
    \wbs_dat_out_3[15] ,
    \wbs_dat_out_3[14] ,
    \wbs_dat_out_3[13] ,
    \wbs_dat_out_3[12] ,
    \wbs_dat_out_3[11] ,
    \wbs_dat_out_3[10] ,
    \wbs_dat_out_3[9] ,
    \wbs_dat_out_3[8] ,
    \wbs_dat_out_3[7] ,
    \wbs_dat_out_3[6] ,
    \wbs_dat_out_3[5] ,
    \wbs_dat_out_3[4] ,
    \wbs_dat_out_3[3] ,
    \wbs_dat_out_3[2] ,
    \wbs_dat_out_3[1] ,
    \wbs_dat_out_3[0] }),
    .m_wbs_dat_o_4({\wbs_dat_out_4[31] ,
    \wbs_dat_out_4[30] ,
    \wbs_dat_out_4[29] ,
    \wbs_dat_out_4[28] ,
    \wbs_dat_out_4[27] ,
    \wbs_dat_out_4[26] ,
    \wbs_dat_out_4[25] ,
    \wbs_dat_out_4[24] ,
    \wbs_dat_out_4[23] ,
    \wbs_dat_out_4[22] ,
    \wbs_dat_out_4[21] ,
    \wbs_dat_out_4[20] ,
    \wbs_dat_out_4[19] ,
    \wbs_dat_out_4[18] ,
    \wbs_dat_out_4[17] ,
    \wbs_dat_out_4[16] ,
    \wbs_dat_out_4[15] ,
    \wbs_dat_out_4[14] ,
    \wbs_dat_out_4[13] ,
    \wbs_dat_out_4[12] ,
    \wbs_dat_out_4[11] ,
    \wbs_dat_out_4[10] ,
    \wbs_dat_out_4[9] ,
    \wbs_dat_out_4[8] ,
    \wbs_dat_out_4[7] ,
    \wbs_dat_out_4[6] ,
    \wbs_dat_out_4[5] ,
    \wbs_dat_out_4[4] ,
    \wbs_dat_out_4[3] ,
    \wbs_dat_out_4[2] ,
    \wbs_dat_out_4[1] ,
    \wbs_dat_out_4[0] }),
    .m_wbs_dat_o_5({\wbs_dat_out_5[31] ,
    \wbs_dat_out_5[30] ,
    \wbs_dat_out_5[29] ,
    \wbs_dat_out_5[28] ,
    \wbs_dat_out_5[27] ,
    \wbs_dat_out_5[26] ,
    \wbs_dat_out_5[25] ,
    \wbs_dat_out_5[24] ,
    \wbs_dat_out_5[23] ,
    \wbs_dat_out_5[22] ,
    \wbs_dat_out_5[21] ,
    \wbs_dat_out_5[20] ,
    \wbs_dat_out_5[19] ,
    \wbs_dat_out_5[18] ,
    \wbs_dat_out_5[17] ,
    \wbs_dat_out_5[16] ,
    \wbs_dat_out_5[15] ,
    \wbs_dat_out_5[14] ,
    \wbs_dat_out_5[13] ,
    \wbs_dat_out_5[12] ,
    \wbs_dat_out_5[11] ,
    \wbs_dat_out_5[10] ,
    \wbs_dat_out_5[9] ,
    \wbs_dat_out_5[8] ,
    \wbs_dat_out_5[7] ,
    \wbs_dat_out_5[6] ,
    \wbs_dat_out_5[5] ,
    \wbs_dat_out_5[4] ,
    \wbs_dat_out_5[3] ,
    \wbs_dat_out_5[2] ,
    \wbs_dat_out_5[1] ,
    \wbs_dat_out_5[0] }),
    .m_wbs_dat_o_6({\wbs_dat_out_6[31] ,
    \wbs_dat_out_6[30] ,
    \wbs_dat_out_6[29] ,
    \wbs_dat_out_6[28] ,
    \wbs_dat_out_6[27] ,
    \wbs_dat_out_6[26] ,
    \wbs_dat_out_6[25] ,
    \wbs_dat_out_6[24] ,
    \wbs_dat_out_6[23] ,
    \wbs_dat_out_6[22] ,
    \wbs_dat_out_6[21] ,
    \wbs_dat_out_6[20] ,
    \wbs_dat_out_6[19] ,
    \wbs_dat_out_6[18] ,
    \wbs_dat_out_6[17] ,
    \wbs_dat_out_6[16] ,
    \wbs_dat_out_6[15] ,
    \wbs_dat_out_6[14] ,
    \wbs_dat_out_6[13] ,
    \wbs_dat_out_6[12] ,
    \wbs_dat_out_6[11] ,
    \wbs_dat_out_6[10] ,
    \wbs_dat_out_6[9] ,
    \wbs_dat_out_6[8] ,
    \wbs_dat_out_6[7] ,
    \wbs_dat_out_6[6] ,
    \wbs_dat_out_6[5] ,
    \wbs_dat_out_6[4] ,
    \wbs_dat_out_6[3] ,
    \wbs_dat_out_6[2] ,
    \wbs_dat_out_6[1] ,
    \wbs_dat_out_6[0] }),
    .m_wbs_dat_o_7({\wbs_dat_out_7[31] ,
    \wbs_dat_out_7[30] ,
    \wbs_dat_out_7[29] ,
    \wbs_dat_out_7[28] ,
    \wbs_dat_out_7[27] ,
    \wbs_dat_out_7[26] ,
    \wbs_dat_out_7[25] ,
    \wbs_dat_out_7[24] ,
    \wbs_dat_out_7[23] ,
    \wbs_dat_out_7[22] ,
    \wbs_dat_out_7[21] ,
    \wbs_dat_out_7[20] ,
    \wbs_dat_out_7[19] ,
    \wbs_dat_out_7[18] ,
    \wbs_dat_out_7[17] ,
    \wbs_dat_out_7[16] ,
    \wbs_dat_out_7[15] ,
    \wbs_dat_out_7[14] ,
    \wbs_dat_out_7[13] ,
    \wbs_dat_out_7[12] ,
    \wbs_dat_out_7[11] ,
    \wbs_dat_out_7[10] ,
    \wbs_dat_out_7[9] ,
    \wbs_dat_out_7[8] ,
    \wbs_dat_out_7[7] ,
    \wbs_dat_out_7[6] ,
    \wbs_dat_out_7[5] ,
    \wbs_dat_out_7[4] ,
    \wbs_dat_out_7[3] ,
    \wbs_dat_out_7[2] ,
    \wbs_dat_out_7[1] ,
    \wbs_dat_out_7[0] }),
    .m_wbs_dat_o_8({\wbs_dat_out_8[31] ,
    \wbs_dat_out_8[30] ,
    \wbs_dat_out_8[29] ,
    \wbs_dat_out_8[28] ,
    \wbs_dat_out_8[27] ,
    \wbs_dat_out_8[26] ,
    \wbs_dat_out_8[25] ,
    \wbs_dat_out_8[24] ,
    \wbs_dat_out_8[23] ,
    \wbs_dat_out_8[22] ,
    \wbs_dat_out_8[21] ,
    \wbs_dat_out_8[20] ,
    \wbs_dat_out_8[19] ,
    \wbs_dat_out_8[18] ,
    \wbs_dat_out_8[17] ,
    \wbs_dat_out_8[16] ,
    \wbs_dat_out_8[15] ,
    \wbs_dat_out_8[14] ,
    \wbs_dat_out_8[13] ,
    \wbs_dat_out_8[12] ,
    \wbs_dat_out_8[11] ,
    \wbs_dat_out_8[10] ,
    \wbs_dat_out_8[9] ,
    \wbs_dat_out_8[8] ,
    \wbs_dat_out_8[7] ,
    \wbs_dat_out_8[6] ,
    \wbs_dat_out_8[5] ,
    \wbs_dat_out_8[4] ,
    \wbs_dat_out_8[3] ,
    \wbs_dat_out_8[2] ,
    \wbs_dat_out_8[1] ,
    \wbs_dat_out_8[0] }),
    .m_wbs_dat_o_9({\wbs_dat_out_9[31] ,
    \wbs_dat_out_9[30] ,
    \wbs_dat_out_9[29] ,
    \wbs_dat_out_9[28] ,
    \wbs_dat_out_9[27] ,
    \wbs_dat_out_9[26] ,
    \wbs_dat_out_9[25] ,
    \wbs_dat_out_9[24] ,
    \wbs_dat_out_9[23] ,
    \wbs_dat_out_9[22] ,
    \wbs_dat_out_9[21] ,
    \wbs_dat_out_9[20] ,
    \wbs_dat_out_9[19] ,
    \wbs_dat_out_9[18] ,
    \wbs_dat_out_9[17] ,
    \wbs_dat_out_9[16] ,
    \wbs_dat_out_9[15] ,
    \wbs_dat_out_9[14] ,
    \wbs_dat_out_9[13] ,
    \wbs_dat_out_9[12] ,
    \wbs_dat_out_9[11] ,
    \wbs_dat_out_9[10] ,
    \wbs_dat_out_9[9] ,
    \wbs_dat_out_9[8] ,
    \wbs_dat_out_9[7] ,
    \wbs_dat_out_9[6] ,
    \wbs_dat_out_9[5] ,
    \wbs_dat_out_9[4] ,
    \wbs_dat_out_9[3] ,
    \wbs_dat_out_9[2] ,
    \wbs_dat_out_9[1] ,
    \wbs_dat_out_9[0] }),
    .m_wbs_stb_i({\m_wbs_stb_i[10] ,
    \m_wbs_stb_i[9] ,
    \m_wbs_stb_i[8] ,
    \m_wbs_stb_i[7] ,
    \m_wbs_stb_i[6] ,
    \m_wbs_stb_i[5] ,
    \m_wbs_stb_i[4] ,
    \m_wbs_stb_i[3] ,
    \m_wbs_stb_i[2] ,
    \m_wbs_stb_i[1] ,
    \m_wbs_stb_i[0] }),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}));
 ren_conv_top ren_conv_top_inst_0 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[0] ),
    .wbs_ack_o(\m_wbs_ack_out[0] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[0] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_0[31] ,
    \wbs_dat_out_0[30] ,
    \wbs_dat_out_0[29] ,
    \wbs_dat_out_0[28] ,
    \wbs_dat_out_0[27] ,
    \wbs_dat_out_0[26] ,
    \wbs_dat_out_0[25] ,
    \wbs_dat_out_0[24] ,
    \wbs_dat_out_0[23] ,
    \wbs_dat_out_0[22] ,
    \wbs_dat_out_0[21] ,
    \wbs_dat_out_0[20] ,
    \wbs_dat_out_0[19] ,
    \wbs_dat_out_0[18] ,
    \wbs_dat_out_0[17] ,
    \wbs_dat_out_0[16] ,
    \wbs_dat_out_0[15] ,
    \wbs_dat_out_0[14] ,
    \wbs_dat_out_0[13] ,
    \wbs_dat_out_0[12] ,
    \wbs_dat_out_0[11] ,
    \wbs_dat_out_0[10] ,
    \wbs_dat_out_0[9] ,
    \wbs_dat_out_0[8] ,
    \wbs_dat_out_0[7] ,
    \wbs_dat_out_0[6] ,
    \wbs_dat_out_0[5] ,
    \wbs_dat_out_0[4] ,
    \wbs_dat_out_0[3] ,
    \wbs_dat_out_0[2] ,
    \wbs_dat_out_0[1] ,
    \wbs_dat_out_0[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_1 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[1] ),
    .wbs_ack_o(\m_wbs_ack_out[1] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[1] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_1[31] ,
    \wbs_dat_out_1[30] ,
    \wbs_dat_out_1[29] ,
    \wbs_dat_out_1[28] ,
    \wbs_dat_out_1[27] ,
    \wbs_dat_out_1[26] ,
    \wbs_dat_out_1[25] ,
    \wbs_dat_out_1[24] ,
    \wbs_dat_out_1[23] ,
    \wbs_dat_out_1[22] ,
    \wbs_dat_out_1[21] ,
    \wbs_dat_out_1[20] ,
    \wbs_dat_out_1[19] ,
    \wbs_dat_out_1[18] ,
    \wbs_dat_out_1[17] ,
    \wbs_dat_out_1[16] ,
    \wbs_dat_out_1[15] ,
    \wbs_dat_out_1[14] ,
    \wbs_dat_out_1[13] ,
    \wbs_dat_out_1[12] ,
    \wbs_dat_out_1[11] ,
    \wbs_dat_out_1[10] ,
    \wbs_dat_out_1[9] ,
    \wbs_dat_out_1[8] ,
    \wbs_dat_out_1[7] ,
    \wbs_dat_out_1[6] ,
    \wbs_dat_out_1[5] ,
    \wbs_dat_out_1[4] ,
    \wbs_dat_out_1[3] ,
    \wbs_dat_out_1[2] ,
    \wbs_dat_out_1[1] ,
    \wbs_dat_out_1[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_10 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[10] ),
    .wbs_ack_o(\m_wbs_ack_out[10] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[10] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_10[31] ,
    \wbs_dat_out_10[30] ,
    \wbs_dat_out_10[29] ,
    \wbs_dat_out_10[28] ,
    \wbs_dat_out_10[27] ,
    \wbs_dat_out_10[26] ,
    \wbs_dat_out_10[25] ,
    \wbs_dat_out_10[24] ,
    \wbs_dat_out_10[23] ,
    \wbs_dat_out_10[22] ,
    \wbs_dat_out_10[21] ,
    \wbs_dat_out_10[20] ,
    \wbs_dat_out_10[19] ,
    \wbs_dat_out_10[18] ,
    \wbs_dat_out_10[17] ,
    \wbs_dat_out_10[16] ,
    \wbs_dat_out_10[15] ,
    \wbs_dat_out_10[14] ,
    \wbs_dat_out_10[13] ,
    \wbs_dat_out_10[12] ,
    \wbs_dat_out_10[11] ,
    \wbs_dat_out_10[10] ,
    \wbs_dat_out_10[9] ,
    \wbs_dat_out_10[8] ,
    \wbs_dat_out_10[7] ,
    \wbs_dat_out_10[6] ,
    \wbs_dat_out_10[5] ,
    \wbs_dat_out_10[4] ,
    \wbs_dat_out_10[3] ,
    \wbs_dat_out_10[2] ,
    \wbs_dat_out_10[1] ,
    \wbs_dat_out_10[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_2 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[2] ),
    .wbs_ack_o(\m_wbs_ack_out[2] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[2] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_2[31] ,
    \wbs_dat_out_2[30] ,
    \wbs_dat_out_2[29] ,
    \wbs_dat_out_2[28] ,
    \wbs_dat_out_2[27] ,
    \wbs_dat_out_2[26] ,
    \wbs_dat_out_2[25] ,
    \wbs_dat_out_2[24] ,
    \wbs_dat_out_2[23] ,
    \wbs_dat_out_2[22] ,
    \wbs_dat_out_2[21] ,
    \wbs_dat_out_2[20] ,
    \wbs_dat_out_2[19] ,
    \wbs_dat_out_2[18] ,
    \wbs_dat_out_2[17] ,
    \wbs_dat_out_2[16] ,
    \wbs_dat_out_2[15] ,
    \wbs_dat_out_2[14] ,
    \wbs_dat_out_2[13] ,
    \wbs_dat_out_2[12] ,
    \wbs_dat_out_2[11] ,
    \wbs_dat_out_2[10] ,
    \wbs_dat_out_2[9] ,
    \wbs_dat_out_2[8] ,
    \wbs_dat_out_2[7] ,
    \wbs_dat_out_2[6] ,
    \wbs_dat_out_2[5] ,
    \wbs_dat_out_2[4] ,
    \wbs_dat_out_2[3] ,
    \wbs_dat_out_2[2] ,
    \wbs_dat_out_2[1] ,
    \wbs_dat_out_2[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_3 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[3] ),
    .wbs_ack_o(\m_wbs_ack_out[3] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[3] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_3[31] ,
    \wbs_dat_out_3[30] ,
    \wbs_dat_out_3[29] ,
    \wbs_dat_out_3[28] ,
    \wbs_dat_out_3[27] ,
    \wbs_dat_out_3[26] ,
    \wbs_dat_out_3[25] ,
    \wbs_dat_out_3[24] ,
    \wbs_dat_out_3[23] ,
    \wbs_dat_out_3[22] ,
    \wbs_dat_out_3[21] ,
    \wbs_dat_out_3[20] ,
    \wbs_dat_out_3[19] ,
    \wbs_dat_out_3[18] ,
    \wbs_dat_out_3[17] ,
    \wbs_dat_out_3[16] ,
    \wbs_dat_out_3[15] ,
    \wbs_dat_out_3[14] ,
    \wbs_dat_out_3[13] ,
    \wbs_dat_out_3[12] ,
    \wbs_dat_out_3[11] ,
    \wbs_dat_out_3[10] ,
    \wbs_dat_out_3[9] ,
    \wbs_dat_out_3[8] ,
    \wbs_dat_out_3[7] ,
    \wbs_dat_out_3[6] ,
    \wbs_dat_out_3[5] ,
    \wbs_dat_out_3[4] ,
    \wbs_dat_out_3[3] ,
    \wbs_dat_out_3[2] ,
    \wbs_dat_out_3[1] ,
    \wbs_dat_out_3[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_4 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[4] ),
    .wbs_ack_o(\m_wbs_ack_out[4] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[4] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_4[31] ,
    \wbs_dat_out_4[30] ,
    \wbs_dat_out_4[29] ,
    \wbs_dat_out_4[28] ,
    \wbs_dat_out_4[27] ,
    \wbs_dat_out_4[26] ,
    \wbs_dat_out_4[25] ,
    \wbs_dat_out_4[24] ,
    \wbs_dat_out_4[23] ,
    \wbs_dat_out_4[22] ,
    \wbs_dat_out_4[21] ,
    \wbs_dat_out_4[20] ,
    \wbs_dat_out_4[19] ,
    \wbs_dat_out_4[18] ,
    \wbs_dat_out_4[17] ,
    \wbs_dat_out_4[16] ,
    \wbs_dat_out_4[15] ,
    \wbs_dat_out_4[14] ,
    \wbs_dat_out_4[13] ,
    \wbs_dat_out_4[12] ,
    \wbs_dat_out_4[11] ,
    \wbs_dat_out_4[10] ,
    \wbs_dat_out_4[9] ,
    \wbs_dat_out_4[8] ,
    \wbs_dat_out_4[7] ,
    \wbs_dat_out_4[6] ,
    \wbs_dat_out_4[5] ,
    \wbs_dat_out_4[4] ,
    \wbs_dat_out_4[3] ,
    \wbs_dat_out_4[2] ,
    \wbs_dat_out_4[1] ,
    \wbs_dat_out_4[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_5 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[5] ),
    .wbs_ack_o(\m_wbs_ack_out[5] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[5] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_5[31] ,
    \wbs_dat_out_5[30] ,
    \wbs_dat_out_5[29] ,
    \wbs_dat_out_5[28] ,
    \wbs_dat_out_5[27] ,
    \wbs_dat_out_5[26] ,
    \wbs_dat_out_5[25] ,
    \wbs_dat_out_5[24] ,
    \wbs_dat_out_5[23] ,
    \wbs_dat_out_5[22] ,
    \wbs_dat_out_5[21] ,
    \wbs_dat_out_5[20] ,
    \wbs_dat_out_5[19] ,
    \wbs_dat_out_5[18] ,
    \wbs_dat_out_5[17] ,
    \wbs_dat_out_5[16] ,
    \wbs_dat_out_5[15] ,
    \wbs_dat_out_5[14] ,
    \wbs_dat_out_5[13] ,
    \wbs_dat_out_5[12] ,
    \wbs_dat_out_5[11] ,
    \wbs_dat_out_5[10] ,
    \wbs_dat_out_5[9] ,
    \wbs_dat_out_5[8] ,
    \wbs_dat_out_5[7] ,
    \wbs_dat_out_5[6] ,
    \wbs_dat_out_5[5] ,
    \wbs_dat_out_5[4] ,
    \wbs_dat_out_5[3] ,
    \wbs_dat_out_5[2] ,
    \wbs_dat_out_5[1] ,
    \wbs_dat_out_5[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_6 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[6] ),
    .wbs_ack_o(\m_wbs_ack_out[6] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[6] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_6[31] ,
    \wbs_dat_out_6[30] ,
    \wbs_dat_out_6[29] ,
    \wbs_dat_out_6[28] ,
    \wbs_dat_out_6[27] ,
    \wbs_dat_out_6[26] ,
    \wbs_dat_out_6[25] ,
    \wbs_dat_out_6[24] ,
    \wbs_dat_out_6[23] ,
    \wbs_dat_out_6[22] ,
    \wbs_dat_out_6[21] ,
    \wbs_dat_out_6[20] ,
    \wbs_dat_out_6[19] ,
    \wbs_dat_out_6[18] ,
    \wbs_dat_out_6[17] ,
    \wbs_dat_out_6[16] ,
    \wbs_dat_out_6[15] ,
    \wbs_dat_out_6[14] ,
    \wbs_dat_out_6[13] ,
    \wbs_dat_out_6[12] ,
    \wbs_dat_out_6[11] ,
    \wbs_dat_out_6[10] ,
    \wbs_dat_out_6[9] ,
    \wbs_dat_out_6[8] ,
    \wbs_dat_out_6[7] ,
    \wbs_dat_out_6[6] ,
    \wbs_dat_out_6[5] ,
    \wbs_dat_out_6[4] ,
    \wbs_dat_out_6[3] ,
    \wbs_dat_out_6[2] ,
    \wbs_dat_out_6[1] ,
    \wbs_dat_out_6[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_7 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[7] ),
    .wbs_ack_o(\m_wbs_ack_out[7] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[7] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_7[31] ,
    \wbs_dat_out_7[30] ,
    \wbs_dat_out_7[29] ,
    \wbs_dat_out_7[28] ,
    \wbs_dat_out_7[27] ,
    \wbs_dat_out_7[26] ,
    \wbs_dat_out_7[25] ,
    \wbs_dat_out_7[24] ,
    \wbs_dat_out_7[23] ,
    \wbs_dat_out_7[22] ,
    \wbs_dat_out_7[21] ,
    \wbs_dat_out_7[20] ,
    \wbs_dat_out_7[19] ,
    \wbs_dat_out_7[18] ,
    \wbs_dat_out_7[17] ,
    \wbs_dat_out_7[16] ,
    \wbs_dat_out_7[15] ,
    \wbs_dat_out_7[14] ,
    \wbs_dat_out_7[13] ,
    \wbs_dat_out_7[12] ,
    \wbs_dat_out_7[11] ,
    \wbs_dat_out_7[10] ,
    \wbs_dat_out_7[9] ,
    \wbs_dat_out_7[8] ,
    \wbs_dat_out_7[7] ,
    \wbs_dat_out_7[6] ,
    \wbs_dat_out_7[5] ,
    \wbs_dat_out_7[4] ,
    \wbs_dat_out_7[3] ,
    \wbs_dat_out_7[2] ,
    \wbs_dat_out_7[1] ,
    \wbs_dat_out_7[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_8 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[8] ),
    .wbs_ack_o(\m_wbs_ack_out[8] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[8] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_8[31] ,
    \wbs_dat_out_8[30] ,
    \wbs_dat_out_8[29] ,
    \wbs_dat_out_8[28] ,
    \wbs_dat_out_8[27] ,
    \wbs_dat_out_8[26] ,
    \wbs_dat_out_8[25] ,
    \wbs_dat_out_8[24] ,
    \wbs_dat_out_8[23] ,
    \wbs_dat_out_8[22] ,
    \wbs_dat_out_8[21] ,
    \wbs_dat_out_8[20] ,
    \wbs_dat_out_8[19] ,
    \wbs_dat_out_8[18] ,
    \wbs_dat_out_8[17] ,
    \wbs_dat_out_8[16] ,
    \wbs_dat_out_8[15] ,
    \wbs_dat_out_8[14] ,
    \wbs_dat_out_8[13] ,
    \wbs_dat_out_8[12] ,
    \wbs_dat_out_8[11] ,
    \wbs_dat_out_8[10] ,
    \wbs_dat_out_8[9] ,
    \wbs_dat_out_8[8] ,
    \wbs_dat_out_8[7] ,
    \wbs_dat_out_8[6] ,
    \wbs_dat_out_8[5] ,
    \wbs_dat_out_8[4] ,
    \wbs_dat_out_8[3] ,
    \wbs_dat_out_8[2] ,
    \wbs_dat_out_8[1] ,
    \wbs_dat_out_8[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
 ren_conv_top ren_conv_top_inst_9 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(\m_wb_rst_i[9] ),
    .wbs_ack_o(\m_wbs_ack_out[9] ),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(\m_wbs_stb_i[9] ),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({\wbs_dat_out_9[31] ,
    \wbs_dat_out_9[30] ,
    \wbs_dat_out_9[29] ,
    \wbs_dat_out_9[28] ,
    \wbs_dat_out_9[27] ,
    \wbs_dat_out_9[26] ,
    \wbs_dat_out_9[25] ,
    \wbs_dat_out_9[24] ,
    \wbs_dat_out_9[23] ,
    \wbs_dat_out_9[22] ,
    \wbs_dat_out_9[21] ,
    \wbs_dat_out_9[20] ,
    \wbs_dat_out_9[19] ,
    \wbs_dat_out_9[18] ,
    \wbs_dat_out_9[17] ,
    \wbs_dat_out_9[16] ,
    \wbs_dat_out_9[15] ,
    \wbs_dat_out_9[14] ,
    \wbs_dat_out_9[13] ,
    \wbs_dat_out_9[12] ,
    \wbs_dat_out_9[11] ,
    \wbs_dat_out_9[10] ,
    \wbs_dat_out_9[9] ,
    \wbs_dat_out_9[8] ,
    \wbs_dat_out_9[7] ,
    \wbs_dat_out_9[6] ,
    \wbs_dat_out_9[5] ,
    \wbs_dat_out_9[4] ,
    \wbs_dat_out_9[3] ,
    \wbs_dat_out_9[2] ,
    \wbs_dat_out_9[1] ,
    \wbs_dat_out_9[0] }),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}));
endmodule
