* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for ren_conv_top abstract view
.subckt ren_conv_top wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for multiplex abstract view
.subckt multiplex io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1]
+ irq[2] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103]
+ la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108]
+ la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112]
+ la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117]
+ la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121]
+ la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126]
+ la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65]
+ la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70]
+ la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75]
+ la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80]
+ la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85]
+ la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90]
+ la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95]
+ la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] m_wb_rst_i[0]
+ m_wb_rst_i[10] m_wb_rst_i[1] m_wb_rst_i[2] m_wb_rst_i[3] m_wb_rst_i[4] m_wb_rst_i[5]
+ m_wb_rst_i[6] m_wb_rst_i[7] m_wb_rst_i[8] m_wb_rst_i[9] m_wbs_ack_o[0] m_wbs_ack_o[10]
+ m_wbs_ack_o[1] m_wbs_ack_o[2] m_wbs_ack_o[3] m_wbs_ack_o[4] m_wbs_ack_o[5] m_wbs_ack_o[6]
+ m_wbs_ack_o[7] m_wbs_ack_o[8] m_wbs_ack_o[9] m_wbs_dat_o_0[0] m_wbs_dat_o_0[10]
+ m_wbs_dat_o_0[11] m_wbs_dat_o_0[12] m_wbs_dat_o_0[13] m_wbs_dat_o_0[14] m_wbs_dat_o_0[15]
+ m_wbs_dat_o_0[16] m_wbs_dat_o_0[17] m_wbs_dat_o_0[18] m_wbs_dat_o_0[19] m_wbs_dat_o_0[1]
+ m_wbs_dat_o_0[20] m_wbs_dat_o_0[21] m_wbs_dat_o_0[22] m_wbs_dat_o_0[23] m_wbs_dat_o_0[24]
+ m_wbs_dat_o_0[25] m_wbs_dat_o_0[26] m_wbs_dat_o_0[27] m_wbs_dat_o_0[28] m_wbs_dat_o_0[29]
+ m_wbs_dat_o_0[2] m_wbs_dat_o_0[30] m_wbs_dat_o_0[31] m_wbs_dat_o_0[3] m_wbs_dat_o_0[4]
+ m_wbs_dat_o_0[5] m_wbs_dat_o_0[6] m_wbs_dat_o_0[7] m_wbs_dat_o_0[8] m_wbs_dat_o_0[9]
+ m_wbs_dat_o_10[0] m_wbs_dat_o_10[10] m_wbs_dat_o_10[11] m_wbs_dat_o_10[12] m_wbs_dat_o_10[13]
+ m_wbs_dat_o_10[14] m_wbs_dat_o_10[15] m_wbs_dat_o_10[16] m_wbs_dat_o_10[17] m_wbs_dat_o_10[18]
+ m_wbs_dat_o_10[19] m_wbs_dat_o_10[1] m_wbs_dat_o_10[20] m_wbs_dat_o_10[21] m_wbs_dat_o_10[22]
+ m_wbs_dat_o_10[23] m_wbs_dat_o_10[24] m_wbs_dat_o_10[25] m_wbs_dat_o_10[26] m_wbs_dat_o_10[27]
+ m_wbs_dat_o_10[28] m_wbs_dat_o_10[29] m_wbs_dat_o_10[2] m_wbs_dat_o_10[30] m_wbs_dat_o_10[31]
+ m_wbs_dat_o_10[3] m_wbs_dat_o_10[4] m_wbs_dat_o_10[5] m_wbs_dat_o_10[6] m_wbs_dat_o_10[7]
+ m_wbs_dat_o_10[8] m_wbs_dat_o_10[9] m_wbs_dat_o_1[0] m_wbs_dat_o_1[10] m_wbs_dat_o_1[11]
+ m_wbs_dat_o_1[12] m_wbs_dat_o_1[13] m_wbs_dat_o_1[14] m_wbs_dat_o_1[15] m_wbs_dat_o_1[16]
+ m_wbs_dat_o_1[17] m_wbs_dat_o_1[18] m_wbs_dat_o_1[19] m_wbs_dat_o_1[1] m_wbs_dat_o_1[20]
+ m_wbs_dat_o_1[21] m_wbs_dat_o_1[22] m_wbs_dat_o_1[23] m_wbs_dat_o_1[24] m_wbs_dat_o_1[25]
+ m_wbs_dat_o_1[26] m_wbs_dat_o_1[27] m_wbs_dat_o_1[28] m_wbs_dat_o_1[29] m_wbs_dat_o_1[2]
+ m_wbs_dat_o_1[30] m_wbs_dat_o_1[31] m_wbs_dat_o_1[3] m_wbs_dat_o_1[4] m_wbs_dat_o_1[5]
+ m_wbs_dat_o_1[6] m_wbs_dat_o_1[7] m_wbs_dat_o_1[8] m_wbs_dat_o_1[9] m_wbs_dat_o_2[0]
+ m_wbs_dat_o_2[10] m_wbs_dat_o_2[11] m_wbs_dat_o_2[12] m_wbs_dat_o_2[13] m_wbs_dat_o_2[14]
+ m_wbs_dat_o_2[15] m_wbs_dat_o_2[16] m_wbs_dat_o_2[17] m_wbs_dat_o_2[18] m_wbs_dat_o_2[19]
+ m_wbs_dat_o_2[1] m_wbs_dat_o_2[20] m_wbs_dat_o_2[21] m_wbs_dat_o_2[22] m_wbs_dat_o_2[23]
+ m_wbs_dat_o_2[24] m_wbs_dat_o_2[25] m_wbs_dat_o_2[26] m_wbs_dat_o_2[27] m_wbs_dat_o_2[28]
+ m_wbs_dat_o_2[29] m_wbs_dat_o_2[2] m_wbs_dat_o_2[30] m_wbs_dat_o_2[31] m_wbs_dat_o_2[3]
+ m_wbs_dat_o_2[4] m_wbs_dat_o_2[5] m_wbs_dat_o_2[6] m_wbs_dat_o_2[7] m_wbs_dat_o_2[8]
+ m_wbs_dat_o_2[9] m_wbs_dat_o_3[0] m_wbs_dat_o_3[10] m_wbs_dat_o_3[11] m_wbs_dat_o_3[12]
+ m_wbs_dat_o_3[13] m_wbs_dat_o_3[14] m_wbs_dat_o_3[15] m_wbs_dat_o_3[16] m_wbs_dat_o_3[17]
+ m_wbs_dat_o_3[18] m_wbs_dat_o_3[19] m_wbs_dat_o_3[1] m_wbs_dat_o_3[20] m_wbs_dat_o_3[21]
+ m_wbs_dat_o_3[22] m_wbs_dat_o_3[23] m_wbs_dat_o_3[24] m_wbs_dat_o_3[25] m_wbs_dat_o_3[26]
+ m_wbs_dat_o_3[27] m_wbs_dat_o_3[28] m_wbs_dat_o_3[29] m_wbs_dat_o_3[2] m_wbs_dat_o_3[30]
+ m_wbs_dat_o_3[31] m_wbs_dat_o_3[3] m_wbs_dat_o_3[4] m_wbs_dat_o_3[5] m_wbs_dat_o_3[6]
+ m_wbs_dat_o_3[7] m_wbs_dat_o_3[8] m_wbs_dat_o_3[9] m_wbs_dat_o_4[0] m_wbs_dat_o_4[10]
+ m_wbs_dat_o_4[11] m_wbs_dat_o_4[12] m_wbs_dat_o_4[13] m_wbs_dat_o_4[14] m_wbs_dat_o_4[15]
+ m_wbs_dat_o_4[16] m_wbs_dat_o_4[17] m_wbs_dat_o_4[18] m_wbs_dat_o_4[19] m_wbs_dat_o_4[1]
+ m_wbs_dat_o_4[20] m_wbs_dat_o_4[21] m_wbs_dat_o_4[22] m_wbs_dat_o_4[23] m_wbs_dat_o_4[24]
+ m_wbs_dat_o_4[25] m_wbs_dat_o_4[26] m_wbs_dat_o_4[27] m_wbs_dat_o_4[28] m_wbs_dat_o_4[29]
+ m_wbs_dat_o_4[2] m_wbs_dat_o_4[30] m_wbs_dat_o_4[31] m_wbs_dat_o_4[3] m_wbs_dat_o_4[4]
+ m_wbs_dat_o_4[5] m_wbs_dat_o_4[6] m_wbs_dat_o_4[7] m_wbs_dat_o_4[8] m_wbs_dat_o_4[9]
+ m_wbs_dat_o_5[0] m_wbs_dat_o_5[10] m_wbs_dat_o_5[11] m_wbs_dat_o_5[12] m_wbs_dat_o_5[13]
+ m_wbs_dat_o_5[14] m_wbs_dat_o_5[15] m_wbs_dat_o_5[16] m_wbs_dat_o_5[17] m_wbs_dat_o_5[18]
+ m_wbs_dat_o_5[19] m_wbs_dat_o_5[1] m_wbs_dat_o_5[20] m_wbs_dat_o_5[21] m_wbs_dat_o_5[22]
+ m_wbs_dat_o_5[23] m_wbs_dat_o_5[24] m_wbs_dat_o_5[25] m_wbs_dat_o_5[26] m_wbs_dat_o_5[27]
+ m_wbs_dat_o_5[28] m_wbs_dat_o_5[29] m_wbs_dat_o_5[2] m_wbs_dat_o_5[30] m_wbs_dat_o_5[31]
+ m_wbs_dat_o_5[3] m_wbs_dat_o_5[4] m_wbs_dat_o_5[5] m_wbs_dat_o_5[6] m_wbs_dat_o_5[7]
+ m_wbs_dat_o_5[8] m_wbs_dat_o_5[9] m_wbs_dat_o_6[0] m_wbs_dat_o_6[10] m_wbs_dat_o_6[11]
+ m_wbs_dat_o_6[12] m_wbs_dat_o_6[13] m_wbs_dat_o_6[14] m_wbs_dat_o_6[15] m_wbs_dat_o_6[16]
+ m_wbs_dat_o_6[17] m_wbs_dat_o_6[18] m_wbs_dat_o_6[19] m_wbs_dat_o_6[1] m_wbs_dat_o_6[20]
+ m_wbs_dat_o_6[21] m_wbs_dat_o_6[22] m_wbs_dat_o_6[23] m_wbs_dat_o_6[24] m_wbs_dat_o_6[25]
+ m_wbs_dat_o_6[26] m_wbs_dat_o_6[27] m_wbs_dat_o_6[28] m_wbs_dat_o_6[29] m_wbs_dat_o_6[2]
+ m_wbs_dat_o_6[30] m_wbs_dat_o_6[31] m_wbs_dat_o_6[3] m_wbs_dat_o_6[4] m_wbs_dat_o_6[5]
+ m_wbs_dat_o_6[6] m_wbs_dat_o_6[7] m_wbs_dat_o_6[8] m_wbs_dat_o_6[9] m_wbs_dat_o_7[0]
+ m_wbs_dat_o_7[10] m_wbs_dat_o_7[11] m_wbs_dat_o_7[12] m_wbs_dat_o_7[13] m_wbs_dat_o_7[14]
+ m_wbs_dat_o_7[15] m_wbs_dat_o_7[16] m_wbs_dat_o_7[17] m_wbs_dat_o_7[18] m_wbs_dat_o_7[19]
+ m_wbs_dat_o_7[1] m_wbs_dat_o_7[20] m_wbs_dat_o_7[21] m_wbs_dat_o_7[22] m_wbs_dat_o_7[23]
+ m_wbs_dat_o_7[24] m_wbs_dat_o_7[25] m_wbs_dat_o_7[26] m_wbs_dat_o_7[27] m_wbs_dat_o_7[28]
+ m_wbs_dat_o_7[29] m_wbs_dat_o_7[2] m_wbs_dat_o_7[30] m_wbs_dat_o_7[31] m_wbs_dat_o_7[3]
+ m_wbs_dat_o_7[4] m_wbs_dat_o_7[5] m_wbs_dat_o_7[6] m_wbs_dat_o_7[7] m_wbs_dat_o_7[8]
+ m_wbs_dat_o_7[9] m_wbs_dat_o_8[0] m_wbs_dat_o_8[10] m_wbs_dat_o_8[11] m_wbs_dat_o_8[12]
+ m_wbs_dat_o_8[13] m_wbs_dat_o_8[14] m_wbs_dat_o_8[15] m_wbs_dat_o_8[16] m_wbs_dat_o_8[17]
+ m_wbs_dat_o_8[18] m_wbs_dat_o_8[19] m_wbs_dat_o_8[1] m_wbs_dat_o_8[20] m_wbs_dat_o_8[21]
+ m_wbs_dat_o_8[22] m_wbs_dat_o_8[23] m_wbs_dat_o_8[24] m_wbs_dat_o_8[25] m_wbs_dat_o_8[26]
+ m_wbs_dat_o_8[27] m_wbs_dat_o_8[28] m_wbs_dat_o_8[29] m_wbs_dat_o_8[2] m_wbs_dat_o_8[30]
+ m_wbs_dat_o_8[31] m_wbs_dat_o_8[3] m_wbs_dat_o_8[4] m_wbs_dat_o_8[5] m_wbs_dat_o_8[6]
+ m_wbs_dat_o_8[7] m_wbs_dat_o_8[8] m_wbs_dat_o_8[9] m_wbs_dat_o_9[0] m_wbs_dat_o_9[10]
+ m_wbs_dat_o_9[11] m_wbs_dat_o_9[12] m_wbs_dat_o_9[13] m_wbs_dat_o_9[14] m_wbs_dat_o_9[15]
+ m_wbs_dat_o_9[16] m_wbs_dat_o_9[17] m_wbs_dat_o_9[18] m_wbs_dat_o_9[19] m_wbs_dat_o_9[1]
+ m_wbs_dat_o_9[20] m_wbs_dat_o_9[21] m_wbs_dat_o_9[22] m_wbs_dat_o_9[23] m_wbs_dat_o_9[24]
+ m_wbs_dat_o_9[25] m_wbs_dat_o_9[26] m_wbs_dat_o_9[27] m_wbs_dat_o_9[28] m_wbs_dat_o_9[29]
+ m_wbs_dat_o_9[2] m_wbs_dat_o_9[30] m_wbs_dat_o_9[31] m_wbs_dat_o_9[3] m_wbs_dat_o_9[4]
+ m_wbs_dat_o_9[5] m_wbs_dat_o_9[6] m_wbs_dat_o_9[7] m_wbs_dat_o_9[8] m_wbs_dat_o_9[9]
+ m_wbs_stb_i[0] m_wbs_stb_i[10] m_wbs_stb_i[1] m_wbs_stb_i[2] m_wbs_stb_i[3] m_wbs_stb_i[4]
+ m_wbs_stb_i[5] m_wbs_stb_i[6] m_wbs_stb_i[7] m_wbs_stb_i[8] m_wbs_stb_i[9] wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i vccd1
+ vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2 vssd2_uq0 vssd2_uq1 vssd2_uq2 vssd2_uq3
+ vssd2_uq4 vssd2_uq5 vssd2_uq6 vssd2_uq7 vssd2_uq8 vssd2_uq9 vssd2_uq10 vssd2_uq11
+ vssd2_uq12 vssd2_uq13 vssd2_uq14 vssd2_uq15 vssd2_uq16 vssd2_uq17 vssd2_uq18 vssd2_uq19
+ vssd2_uq20 vssd2_uq21 vdda2_uq0 vdda2_uq1 vdda2_uq2 vdda2_uq3 vdda2_uq4 vdda2_uq5
+ vdda2_uq6 vdda2_uq7 vdda2_uq8 vdda2_uq9 vdda2_uq10 vdda2_uq11 vdda2_uq12 vdda2_uq13
+ vdda2_uq14 vdda2_uq15 vdda2_uq16 vdda2_uq17 vdda2_uq18 vdda2_uq19 vdda2_uq20 vdda2_uq21
+ vdda2_uq22 vdda2_uq23 vdda2_uq24 vdda2_uq25 vdda1_uq0 vdda1_uq1 vdda1_uq2 vdda1_uq3
+ vdda1_uq4 vdda1_uq5 vdda1_uq6 vdda1_uq7 vdda1_uq8 vdda1_uq9 vdda1_uq10 vdda1_uq11
+ vdda1_uq12 vdda1_uq13 vdda1_uq14 vdda1_uq15 vdda1_uq16 vdda1_uq17 vdda1_uq18 vdda1_uq19
+ vdda1_uq20 vdda1_uq21 vdda1_uq22 vdda1_uq23 vccd2_uq0 vccd2_uq1 vccd2_uq2 vccd2_uq3
+ vccd2_uq4 vccd2_uq5 vccd2_uq6 vccd2_uq7 vccd2_uq8 vccd2_uq9 vccd2_uq10 vccd2_uq11
+ vccd2_uq12 vccd2_uq13 vccd2_uq14 vccd2_uq15 vccd2_uq16 vccd2_uq17 vccd2_uq18 vccd2_uq19
+ vccd2_uq20 vccd2_uq21 vccd2_uq22 vccd2_uq23 vccd2_uq24 vccd2_uq25 vssa2_uq0 vssa2_uq1
+ vssa2_uq2 vssa2_uq3 vssa2_uq4 vssa2_uq5 vssa2_uq6 vssa2_uq7 vssa2_uq8 vssa2_uq9
+ vssa2_uq10 vssa2_uq11 vssa2_uq12 vssa2_uq13 vssa2_uq14 vssa2_uq15 vssa2_uq16 vssa2_uq17
+ vssa2_uq18 vssa2_uq19 vssa2_uq20 vssa2_uq21 vssa1_uq0 vssa1_uq1 vssa1_uq2 vssa1_uq3
+ vssa1_uq4 vssa1_uq5 vssa1_uq6 vssa1_uq7 vssa1_uq8
Xren_conv_top_inst_10 wb_clk_i icon/m_wb_rst_i[10] icon/m_wbs_ack_o[10] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_10[0] icon/m_wbs_dat_o_10[10] icon/m_wbs_dat_o_10[11]
+ icon/m_wbs_dat_o_10[12] icon/m_wbs_dat_o_10[13] icon/m_wbs_dat_o_10[14] icon/m_wbs_dat_o_10[15]
+ icon/m_wbs_dat_o_10[16] icon/m_wbs_dat_o_10[17] icon/m_wbs_dat_o_10[18] icon/m_wbs_dat_o_10[19]
+ icon/m_wbs_dat_o_10[1] icon/m_wbs_dat_o_10[20] icon/m_wbs_dat_o_10[21] icon/m_wbs_dat_o_10[22]
+ icon/m_wbs_dat_o_10[23] icon/m_wbs_dat_o_10[24] icon/m_wbs_dat_o_10[25] icon/m_wbs_dat_o_10[26]
+ icon/m_wbs_dat_o_10[27] icon/m_wbs_dat_o_10[28] icon/m_wbs_dat_o_10[29] icon/m_wbs_dat_o_10[2]
+ icon/m_wbs_dat_o_10[30] icon/m_wbs_dat_o_10[31] icon/m_wbs_dat_o_10[3] icon/m_wbs_dat_o_10[4]
+ icon/m_wbs_dat_o_10[5] icon/m_wbs_dat_o_10[6] icon/m_wbs_dat_o_10[7] icon/m_wbs_dat_o_10[8]
+ icon/m_wbs_dat_o_10[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[10]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_0 wb_clk_i icon/m_wb_rst_i[0] icon/m_wbs_ack_o[0] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_0[0] icon/m_wbs_dat_o_0[10] icon/m_wbs_dat_o_0[11]
+ icon/m_wbs_dat_o_0[12] icon/m_wbs_dat_o_0[13] icon/m_wbs_dat_o_0[14] icon/m_wbs_dat_o_0[15]
+ icon/m_wbs_dat_o_0[16] icon/m_wbs_dat_o_0[17] icon/m_wbs_dat_o_0[18] icon/m_wbs_dat_o_0[19]
+ icon/m_wbs_dat_o_0[1] icon/m_wbs_dat_o_0[20] icon/m_wbs_dat_o_0[21] icon/m_wbs_dat_o_0[22]
+ icon/m_wbs_dat_o_0[23] icon/m_wbs_dat_o_0[24] icon/m_wbs_dat_o_0[25] icon/m_wbs_dat_o_0[26]
+ icon/m_wbs_dat_o_0[27] icon/m_wbs_dat_o_0[28] icon/m_wbs_dat_o_0[29] icon/m_wbs_dat_o_0[2]
+ icon/m_wbs_dat_o_0[30] icon/m_wbs_dat_o_0[31] icon/m_wbs_dat_o_0[3] icon/m_wbs_dat_o_0[4]
+ icon/m_wbs_dat_o_0[5] icon/m_wbs_dat_o_0[6] icon/m_wbs_dat_o_0[7] icon/m_wbs_dat_o_0[8]
+ icon/m_wbs_dat_o_0[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[0]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_1 wb_clk_i icon/m_wb_rst_i[1] icon/m_wbs_ack_o[1] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_1[0] icon/m_wbs_dat_o_1[10] icon/m_wbs_dat_o_1[11]
+ icon/m_wbs_dat_o_1[12] icon/m_wbs_dat_o_1[13] icon/m_wbs_dat_o_1[14] icon/m_wbs_dat_o_1[15]
+ icon/m_wbs_dat_o_1[16] icon/m_wbs_dat_o_1[17] icon/m_wbs_dat_o_1[18] icon/m_wbs_dat_o_1[19]
+ icon/m_wbs_dat_o_1[1] icon/m_wbs_dat_o_1[20] icon/m_wbs_dat_o_1[21] icon/m_wbs_dat_o_1[22]
+ icon/m_wbs_dat_o_1[23] icon/m_wbs_dat_o_1[24] icon/m_wbs_dat_o_1[25] icon/m_wbs_dat_o_1[26]
+ icon/m_wbs_dat_o_1[27] icon/m_wbs_dat_o_1[28] icon/m_wbs_dat_o_1[29] icon/m_wbs_dat_o_1[2]
+ icon/m_wbs_dat_o_1[30] icon/m_wbs_dat_o_1[31] icon/m_wbs_dat_o_1[3] icon/m_wbs_dat_o_1[4]
+ icon/m_wbs_dat_o_1[5] icon/m_wbs_dat_o_1[6] icon/m_wbs_dat_o_1[7] icon/m_wbs_dat_o_1[8]
+ icon/m_wbs_dat_o_1[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[1]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_2 wb_clk_i icon/m_wb_rst_i[2] icon/m_wbs_ack_o[2] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_2[0] icon/m_wbs_dat_o_2[10] icon/m_wbs_dat_o_2[11]
+ icon/m_wbs_dat_o_2[12] icon/m_wbs_dat_o_2[13] icon/m_wbs_dat_o_2[14] icon/m_wbs_dat_o_2[15]
+ icon/m_wbs_dat_o_2[16] icon/m_wbs_dat_o_2[17] icon/m_wbs_dat_o_2[18] icon/m_wbs_dat_o_2[19]
+ icon/m_wbs_dat_o_2[1] icon/m_wbs_dat_o_2[20] icon/m_wbs_dat_o_2[21] icon/m_wbs_dat_o_2[22]
+ icon/m_wbs_dat_o_2[23] icon/m_wbs_dat_o_2[24] icon/m_wbs_dat_o_2[25] icon/m_wbs_dat_o_2[26]
+ icon/m_wbs_dat_o_2[27] icon/m_wbs_dat_o_2[28] icon/m_wbs_dat_o_2[29] icon/m_wbs_dat_o_2[2]
+ icon/m_wbs_dat_o_2[30] icon/m_wbs_dat_o_2[31] icon/m_wbs_dat_o_2[3] icon/m_wbs_dat_o_2[4]
+ icon/m_wbs_dat_o_2[5] icon/m_wbs_dat_o_2[6] icon/m_wbs_dat_o_2[7] icon/m_wbs_dat_o_2[8]
+ icon/m_wbs_dat_o_2[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[2]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_3 wb_clk_i icon/m_wb_rst_i[3] icon/m_wbs_ack_o[3] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_3[0] icon/m_wbs_dat_o_3[10] icon/m_wbs_dat_o_3[11]
+ icon/m_wbs_dat_o_3[12] icon/m_wbs_dat_o_3[13] icon/m_wbs_dat_o_3[14] icon/m_wbs_dat_o_3[15]
+ icon/m_wbs_dat_o_3[16] icon/m_wbs_dat_o_3[17] icon/m_wbs_dat_o_3[18] icon/m_wbs_dat_o_3[19]
+ icon/m_wbs_dat_o_3[1] icon/m_wbs_dat_o_3[20] icon/m_wbs_dat_o_3[21] icon/m_wbs_dat_o_3[22]
+ icon/m_wbs_dat_o_3[23] icon/m_wbs_dat_o_3[24] icon/m_wbs_dat_o_3[25] icon/m_wbs_dat_o_3[26]
+ icon/m_wbs_dat_o_3[27] icon/m_wbs_dat_o_3[28] icon/m_wbs_dat_o_3[29] icon/m_wbs_dat_o_3[2]
+ icon/m_wbs_dat_o_3[30] icon/m_wbs_dat_o_3[31] icon/m_wbs_dat_o_3[3] icon/m_wbs_dat_o_3[4]
+ icon/m_wbs_dat_o_3[5] icon/m_wbs_dat_o_3[6] icon/m_wbs_dat_o_3[7] icon/m_wbs_dat_o_3[8]
+ icon/m_wbs_dat_o_3[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[3]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_4 wb_clk_i icon/m_wb_rst_i[4] icon/m_wbs_ack_o[4] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_4[0] icon/m_wbs_dat_o_4[10] icon/m_wbs_dat_o_4[11]
+ icon/m_wbs_dat_o_4[12] icon/m_wbs_dat_o_4[13] icon/m_wbs_dat_o_4[14] icon/m_wbs_dat_o_4[15]
+ icon/m_wbs_dat_o_4[16] icon/m_wbs_dat_o_4[17] icon/m_wbs_dat_o_4[18] icon/m_wbs_dat_o_4[19]
+ icon/m_wbs_dat_o_4[1] icon/m_wbs_dat_o_4[20] icon/m_wbs_dat_o_4[21] icon/m_wbs_dat_o_4[22]
+ icon/m_wbs_dat_o_4[23] icon/m_wbs_dat_o_4[24] icon/m_wbs_dat_o_4[25] icon/m_wbs_dat_o_4[26]
+ icon/m_wbs_dat_o_4[27] icon/m_wbs_dat_o_4[28] icon/m_wbs_dat_o_4[29] icon/m_wbs_dat_o_4[2]
+ icon/m_wbs_dat_o_4[30] icon/m_wbs_dat_o_4[31] icon/m_wbs_dat_o_4[3] icon/m_wbs_dat_o_4[4]
+ icon/m_wbs_dat_o_4[5] icon/m_wbs_dat_o_4[6] icon/m_wbs_dat_o_4[7] icon/m_wbs_dat_o_4[8]
+ icon/m_wbs_dat_o_4[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[4]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_5 wb_clk_i icon/m_wb_rst_i[5] icon/m_wbs_ack_o[5] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_5[0] icon/m_wbs_dat_o_5[10] icon/m_wbs_dat_o_5[11]
+ icon/m_wbs_dat_o_5[12] icon/m_wbs_dat_o_5[13] icon/m_wbs_dat_o_5[14] icon/m_wbs_dat_o_5[15]
+ icon/m_wbs_dat_o_5[16] icon/m_wbs_dat_o_5[17] icon/m_wbs_dat_o_5[18] icon/m_wbs_dat_o_5[19]
+ icon/m_wbs_dat_o_5[1] icon/m_wbs_dat_o_5[20] icon/m_wbs_dat_o_5[21] icon/m_wbs_dat_o_5[22]
+ icon/m_wbs_dat_o_5[23] icon/m_wbs_dat_o_5[24] icon/m_wbs_dat_o_5[25] icon/m_wbs_dat_o_5[26]
+ icon/m_wbs_dat_o_5[27] icon/m_wbs_dat_o_5[28] icon/m_wbs_dat_o_5[29] icon/m_wbs_dat_o_5[2]
+ icon/m_wbs_dat_o_5[30] icon/m_wbs_dat_o_5[31] icon/m_wbs_dat_o_5[3] icon/m_wbs_dat_o_5[4]
+ icon/m_wbs_dat_o_5[5] icon/m_wbs_dat_o_5[6] icon/m_wbs_dat_o_5[7] icon/m_wbs_dat_o_5[8]
+ icon/m_wbs_dat_o_5[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[5]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_6 wb_clk_i icon/m_wb_rst_i[6] icon/m_wbs_ack_o[6] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_6[0] icon/m_wbs_dat_o_6[10] icon/m_wbs_dat_o_6[11]
+ icon/m_wbs_dat_o_6[12] icon/m_wbs_dat_o_6[13] icon/m_wbs_dat_o_6[14] icon/m_wbs_dat_o_6[15]
+ icon/m_wbs_dat_o_6[16] icon/m_wbs_dat_o_6[17] icon/m_wbs_dat_o_6[18] icon/m_wbs_dat_o_6[19]
+ icon/m_wbs_dat_o_6[1] icon/m_wbs_dat_o_6[20] icon/m_wbs_dat_o_6[21] icon/m_wbs_dat_o_6[22]
+ icon/m_wbs_dat_o_6[23] icon/m_wbs_dat_o_6[24] icon/m_wbs_dat_o_6[25] icon/m_wbs_dat_o_6[26]
+ icon/m_wbs_dat_o_6[27] icon/m_wbs_dat_o_6[28] icon/m_wbs_dat_o_6[29] icon/m_wbs_dat_o_6[2]
+ icon/m_wbs_dat_o_6[30] icon/m_wbs_dat_o_6[31] icon/m_wbs_dat_o_6[3] icon/m_wbs_dat_o_6[4]
+ icon/m_wbs_dat_o_6[5] icon/m_wbs_dat_o_6[6] icon/m_wbs_dat_o_6[7] icon/m_wbs_dat_o_6[8]
+ icon/m_wbs_dat_o_6[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[6]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xicon io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16]
+ io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24]
+ io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32]
+ io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] user_irq[0]
+ user_irq[1] user_irq[2] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] icon/m_wb_rst_i[0] icon/m_wb_rst_i[10] icon/m_wb_rst_i[1] icon/m_wb_rst_i[2]
+ icon/m_wb_rst_i[3] icon/m_wb_rst_i[4] icon/m_wb_rst_i[5] icon/m_wb_rst_i[6] icon/m_wb_rst_i[7]
+ icon/m_wb_rst_i[8] icon/m_wb_rst_i[9] icon/m_wbs_ack_o[0] icon/m_wbs_ack_o[10] icon/m_wbs_ack_o[1]
+ icon/m_wbs_ack_o[2] icon/m_wbs_ack_o[3] icon/m_wbs_ack_o[4] icon/m_wbs_ack_o[5]
+ icon/m_wbs_ack_o[6] icon/m_wbs_ack_o[7] icon/m_wbs_ack_o[8] icon/m_wbs_ack_o[9]
+ icon/m_wbs_dat_o_0[0] icon/m_wbs_dat_o_0[10] icon/m_wbs_dat_o_0[11] icon/m_wbs_dat_o_0[12]
+ icon/m_wbs_dat_o_0[13] icon/m_wbs_dat_o_0[14] icon/m_wbs_dat_o_0[15] icon/m_wbs_dat_o_0[16]
+ icon/m_wbs_dat_o_0[17] icon/m_wbs_dat_o_0[18] icon/m_wbs_dat_o_0[19] icon/m_wbs_dat_o_0[1]
+ icon/m_wbs_dat_o_0[20] icon/m_wbs_dat_o_0[21] icon/m_wbs_dat_o_0[22] icon/m_wbs_dat_o_0[23]
+ icon/m_wbs_dat_o_0[24] icon/m_wbs_dat_o_0[25] icon/m_wbs_dat_o_0[26] icon/m_wbs_dat_o_0[27]
+ icon/m_wbs_dat_o_0[28] icon/m_wbs_dat_o_0[29] icon/m_wbs_dat_o_0[2] icon/m_wbs_dat_o_0[30]
+ icon/m_wbs_dat_o_0[31] icon/m_wbs_dat_o_0[3] icon/m_wbs_dat_o_0[4] icon/m_wbs_dat_o_0[5]
+ icon/m_wbs_dat_o_0[6] icon/m_wbs_dat_o_0[7] icon/m_wbs_dat_o_0[8] icon/m_wbs_dat_o_0[9]
+ icon/m_wbs_dat_o_10[0] icon/m_wbs_dat_o_10[10] icon/m_wbs_dat_o_10[11] icon/m_wbs_dat_o_10[12]
+ icon/m_wbs_dat_o_10[13] icon/m_wbs_dat_o_10[14] icon/m_wbs_dat_o_10[15] icon/m_wbs_dat_o_10[16]
+ icon/m_wbs_dat_o_10[17] icon/m_wbs_dat_o_10[18] icon/m_wbs_dat_o_10[19] icon/m_wbs_dat_o_10[1]
+ icon/m_wbs_dat_o_10[20] icon/m_wbs_dat_o_10[21] icon/m_wbs_dat_o_10[22] icon/m_wbs_dat_o_10[23]
+ icon/m_wbs_dat_o_10[24] icon/m_wbs_dat_o_10[25] icon/m_wbs_dat_o_10[26] icon/m_wbs_dat_o_10[27]
+ icon/m_wbs_dat_o_10[28] icon/m_wbs_dat_o_10[29] icon/m_wbs_dat_o_10[2] icon/m_wbs_dat_o_10[30]
+ icon/m_wbs_dat_o_10[31] icon/m_wbs_dat_o_10[3] icon/m_wbs_dat_o_10[4] icon/m_wbs_dat_o_10[5]
+ icon/m_wbs_dat_o_10[6] icon/m_wbs_dat_o_10[7] icon/m_wbs_dat_o_10[8] icon/m_wbs_dat_o_10[9]
+ icon/m_wbs_dat_o_1[0] icon/m_wbs_dat_o_1[10] icon/m_wbs_dat_o_1[11] icon/m_wbs_dat_o_1[12]
+ icon/m_wbs_dat_o_1[13] icon/m_wbs_dat_o_1[14] icon/m_wbs_dat_o_1[15] icon/m_wbs_dat_o_1[16]
+ icon/m_wbs_dat_o_1[17] icon/m_wbs_dat_o_1[18] icon/m_wbs_dat_o_1[19] icon/m_wbs_dat_o_1[1]
+ icon/m_wbs_dat_o_1[20] icon/m_wbs_dat_o_1[21] icon/m_wbs_dat_o_1[22] icon/m_wbs_dat_o_1[23]
+ icon/m_wbs_dat_o_1[24] icon/m_wbs_dat_o_1[25] icon/m_wbs_dat_o_1[26] icon/m_wbs_dat_o_1[27]
+ icon/m_wbs_dat_o_1[28] icon/m_wbs_dat_o_1[29] icon/m_wbs_dat_o_1[2] icon/m_wbs_dat_o_1[30]
+ icon/m_wbs_dat_o_1[31] icon/m_wbs_dat_o_1[3] icon/m_wbs_dat_o_1[4] icon/m_wbs_dat_o_1[5]
+ icon/m_wbs_dat_o_1[6] icon/m_wbs_dat_o_1[7] icon/m_wbs_dat_o_1[8] icon/m_wbs_dat_o_1[9]
+ icon/m_wbs_dat_o_2[0] icon/m_wbs_dat_o_2[10] icon/m_wbs_dat_o_2[11] icon/m_wbs_dat_o_2[12]
+ icon/m_wbs_dat_o_2[13] icon/m_wbs_dat_o_2[14] icon/m_wbs_dat_o_2[15] icon/m_wbs_dat_o_2[16]
+ icon/m_wbs_dat_o_2[17] icon/m_wbs_dat_o_2[18] icon/m_wbs_dat_o_2[19] icon/m_wbs_dat_o_2[1]
+ icon/m_wbs_dat_o_2[20] icon/m_wbs_dat_o_2[21] icon/m_wbs_dat_o_2[22] icon/m_wbs_dat_o_2[23]
+ icon/m_wbs_dat_o_2[24] icon/m_wbs_dat_o_2[25] icon/m_wbs_dat_o_2[26] icon/m_wbs_dat_o_2[27]
+ icon/m_wbs_dat_o_2[28] icon/m_wbs_dat_o_2[29] icon/m_wbs_dat_o_2[2] icon/m_wbs_dat_o_2[30]
+ icon/m_wbs_dat_o_2[31] icon/m_wbs_dat_o_2[3] icon/m_wbs_dat_o_2[4] icon/m_wbs_dat_o_2[5]
+ icon/m_wbs_dat_o_2[6] icon/m_wbs_dat_o_2[7] icon/m_wbs_dat_o_2[8] icon/m_wbs_dat_o_2[9]
+ icon/m_wbs_dat_o_3[0] icon/m_wbs_dat_o_3[10] icon/m_wbs_dat_o_3[11] icon/m_wbs_dat_o_3[12]
+ icon/m_wbs_dat_o_3[13] icon/m_wbs_dat_o_3[14] icon/m_wbs_dat_o_3[15] icon/m_wbs_dat_o_3[16]
+ icon/m_wbs_dat_o_3[17] icon/m_wbs_dat_o_3[18] icon/m_wbs_dat_o_3[19] icon/m_wbs_dat_o_3[1]
+ icon/m_wbs_dat_o_3[20] icon/m_wbs_dat_o_3[21] icon/m_wbs_dat_o_3[22] icon/m_wbs_dat_o_3[23]
+ icon/m_wbs_dat_o_3[24] icon/m_wbs_dat_o_3[25] icon/m_wbs_dat_o_3[26] icon/m_wbs_dat_o_3[27]
+ icon/m_wbs_dat_o_3[28] icon/m_wbs_dat_o_3[29] icon/m_wbs_dat_o_3[2] icon/m_wbs_dat_o_3[30]
+ icon/m_wbs_dat_o_3[31] icon/m_wbs_dat_o_3[3] icon/m_wbs_dat_o_3[4] icon/m_wbs_dat_o_3[5]
+ icon/m_wbs_dat_o_3[6] icon/m_wbs_dat_o_3[7] icon/m_wbs_dat_o_3[8] icon/m_wbs_dat_o_3[9]
+ icon/m_wbs_dat_o_4[0] icon/m_wbs_dat_o_4[10] icon/m_wbs_dat_o_4[11] icon/m_wbs_dat_o_4[12]
+ icon/m_wbs_dat_o_4[13] icon/m_wbs_dat_o_4[14] icon/m_wbs_dat_o_4[15] icon/m_wbs_dat_o_4[16]
+ icon/m_wbs_dat_o_4[17] icon/m_wbs_dat_o_4[18] icon/m_wbs_dat_o_4[19] icon/m_wbs_dat_o_4[1]
+ icon/m_wbs_dat_o_4[20] icon/m_wbs_dat_o_4[21] icon/m_wbs_dat_o_4[22] icon/m_wbs_dat_o_4[23]
+ icon/m_wbs_dat_o_4[24] icon/m_wbs_dat_o_4[25] icon/m_wbs_dat_o_4[26] icon/m_wbs_dat_o_4[27]
+ icon/m_wbs_dat_o_4[28] icon/m_wbs_dat_o_4[29] icon/m_wbs_dat_o_4[2] icon/m_wbs_dat_o_4[30]
+ icon/m_wbs_dat_o_4[31] icon/m_wbs_dat_o_4[3] icon/m_wbs_dat_o_4[4] icon/m_wbs_dat_o_4[5]
+ icon/m_wbs_dat_o_4[6] icon/m_wbs_dat_o_4[7] icon/m_wbs_dat_o_4[8] icon/m_wbs_dat_o_4[9]
+ icon/m_wbs_dat_o_5[0] icon/m_wbs_dat_o_5[10] icon/m_wbs_dat_o_5[11] icon/m_wbs_dat_o_5[12]
+ icon/m_wbs_dat_o_5[13] icon/m_wbs_dat_o_5[14] icon/m_wbs_dat_o_5[15] icon/m_wbs_dat_o_5[16]
+ icon/m_wbs_dat_o_5[17] icon/m_wbs_dat_o_5[18] icon/m_wbs_dat_o_5[19] icon/m_wbs_dat_o_5[1]
+ icon/m_wbs_dat_o_5[20] icon/m_wbs_dat_o_5[21] icon/m_wbs_dat_o_5[22] icon/m_wbs_dat_o_5[23]
+ icon/m_wbs_dat_o_5[24] icon/m_wbs_dat_o_5[25] icon/m_wbs_dat_o_5[26] icon/m_wbs_dat_o_5[27]
+ icon/m_wbs_dat_o_5[28] icon/m_wbs_dat_o_5[29] icon/m_wbs_dat_o_5[2] icon/m_wbs_dat_o_5[30]
+ icon/m_wbs_dat_o_5[31] icon/m_wbs_dat_o_5[3] icon/m_wbs_dat_o_5[4] icon/m_wbs_dat_o_5[5]
+ icon/m_wbs_dat_o_5[6] icon/m_wbs_dat_o_5[7] icon/m_wbs_dat_o_5[8] icon/m_wbs_dat_o_5[9]
+ icon/m_wbs_dat_o_6[0] icon/m_wbs_dat_o_6[10] icon/m_wbs_dat_o_6[11] icon/m_wbs_dat_o_6[12]
+ icon/m_wbs_dat_o_6[13] icon/m_wbs_dat_o_6[14] icon/m_wbs_dat_o_6[15] icon/m_wbs_dat_o_6[16]
+ icon/m_wbs_dat_o_6[17] icon/m_wbs_dat_o_6[18] icon/m_wbs_dat_o_6[19] icon/m_wbs_dat_o_6[1]
+ icon/m_wbs_dat_o_6[20] icon/m_wbs_dat_o_6[21] icon/m_wbs_dat_o_6[22] icon/m_wbs_dat_o_6[23]
+ icon/m_wbs_dat_o_6[24] icon/m_wbs_dat_o_6[25] icon/m_wbs_dat_o_6[26] icon/m_wbs_dat_o_6[27]
+ icon/m_wbs_dat_o_6[28] icon/m_wbs_dat_o_6[29] icon/m_wbs_dat_o_6[2] icon/m_wbs_dat_o_6[30]
+ icon/m_wbs_dat_o_6[31] icon/m_wbs_dat_o_6[3] icon/m_wbs_dat_o_6[4] icon/m_wbs_dat_o_6[5]
+ icon/m_wbs_dat_o_6[6] icon/m_wbs_dat_o_6[7] icon/m_wbs_dat_o_6[8] icon/m_wbs_dat_o_6[9]
+ icon/m_wbs_dat_o_7[0] icon/m_wbs_dat_o_7[10] icon/m_wbs_dat_o_7[11] icon/m_wbs_dat_o_7[12]
+ icon/m_wbs_dat_o_7[13] icon/m_wbs_dat_o_7[14] icon/m_wbs_dat_o_7[15] icon/m_wbs_dat_o_7[16]
+ icon/m_wbs_dat_o_7[17] icon/m_wbs_dat_o_7[18] icon/m_wbs_dat_o_7[19] icon/m_wbs_dat_o_7[1]
+ icon/m_wbs_dat_o_7[20] icon/m_wbs_dat_o_7[21] icon/m_wbs_dat_o_7[22] icon/m_wbs_dat_o_7[23]
+ icon/m_wbs_dat_o_7[24] icon/m_wbs_dat_o_7[25] icon/m_wbs_dat_o_7[26] icon/m_wbs_dat_o_7[27]
+ icon/m_wbs_dat_o_7[28] icon/m_wbs_dat_o_7[29] icon/m_wbs_dat_o_7[2] icon/m_wbs_dat_o_7[30]
+ icon/m_wbs_dat_o_7[31] icon/m_wbs_dat_o_7[3] icon/m_wbs_dat_o_7[4] icon/m_wbs_dat_o_7[5]
+ icon/m_wbs_dat_o_7[6] icon/m_wbs_dat_o_7[7] icon/m_wbs_dat_o_7[8] icon/m_wbs_dat_o_7[9]
+ icon/m_wbs_dat_o_8[0] icon/m_wbs_dat_o_8[10] icon/m_wbs_dat_o_8[11] icon/m_wbs_dat_o_8[12]
+ icon/m_wbs_dat_o_8[13] icon/m_wbs_dat_o_8[14] icon/m_wbs_dat_o_8[15] icon/m_wbs_dat_o_8[16]
+ icon/m_wbs_dat_o_8[17] icon/m_wbs_dat_o_8[18] icon/m_wbs_dat_o_8[19] icon/m_wbs_dat_o_8[1]
+ icon/m_wbs_dat_o_8[20] icon/m_wbs_dat_o_8[21] icon/m_wbs_dat_o_8[22] icon/m_wbs_dat_o_8[23]
+ icon/m_wbs_dat_o_8[24] icon/m_wbs_dat_o_8[25] icon/m_wbs_dat_o_8[26] icon/m_wbs_dat_o_8[27]
+ icon/m_wbs_dat_o_8[28] icon/m_wbs_dat_o_8[29] icon/m_wbs_dat_o_8[2] icon/m_wbs_dat_o_8[30]
+ icon/m_wbs_dat_o_8[31] icon/m_wbs_dat_o_8[3] icon/m_wbs_dat_o_8[4] icon/m_wbs_dat_o_8[5]
+ icon/m_wbs_dat_o_8[6] icon/m_wbs_dat_o_8[7] icon/m_wbs_dat_o_8[8] icon/m_wbs_dat_o_8[9]
+ icon/m_wbs_dat_o_9[0] icon/m_wbs_dat_o_9[10] icon/m_wbs_dat_o_9[11] icon/m_wbs_dat_o_9[12]
+ icon/m_wbs_dat_o_9[13] icon/m_wbs_dat_o_9[14] icon/m_wbs_dat_o_9[15] icon/m_wbs_dat_o_9[16]
+ icon/m_wbs_dat_o_9[17] icon/m_wbs_dat_o_9[18] icon/m_wbs_dat_o_9[19] icon/m_wbs_dat_o_9[1]
+ icon/m_wbs_dat_o_9[20] icon/m_wbs_dat_o_9[21] icon/m_wbs_dat_o_9[22] icon/m_wbs_dat_o_9[23]
+ icon/m_wbs_dat_o_9[24] icon/m_wbs_dat_o_9[25] icon/m_wbs_dat_o_9[26] icon/m_wbs_dat_o_9[27]
+ icon/m_wbs_dat_o_9[28] icon/m_wbs_dat_o_9[29] icon/m_wbs_dat_o_9[2] icon/m_wbs_dat_o_9[30]
+ icon/m_wbs_dat_o_9[31] icon/m_wbs_dat_o_9[3] icon/m_wbs_dat_o_9[4] icon/m_wbs_dat_o_9[5]
+ icon/m_wbs_dat_o_9[6] icon/m_wbs_dat_o_9[7] icon/m_wbs_dat_o_9[8] icon/m_wbs_dat_o_9[9]
+ icon/m_wbs_stb_i[0] icon/m_wbs_stb_i[10] icon/m_wbs_stb_i[1] icon/m_wbs_stb_i[2]
+ icon/m_wbs_stb_i[3] icon/m_wbs_stb_i[4] icon/m_wbs_stb_i[5] icon/m_wbs_stb_i[6]
+ icon/m_wbs_stb_i[7] icon/m_wbs_stb_i[8] icon/m_wbs_stb_i[9] wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i vccd1 vssd1 multiplex
Xren_conv_top_inst_8 wb_clk_i icon/m_wb_rst_i[8] icon/m_wbs_ack_o[8] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_8[0] icon/m_wbs_dat_o_8[10] icon/m_wbs_dat_o_8[11]
+ icon/m_wbs_dat_o_8[12] icon/m_wbs_dat_o_8[13] icon/m_wbs_dat_o_8[14] icon/m_wbs_dat_o_8[15]
+ icon/m_wbs_dat_o_8[16] icon/m_wbs_dat_o_8[17] icon/m_wbs_dat_o_8[18] icon/m_wbs_dat_o_8[19]
+ icon/m_wbs_dat_o_8[1] icon/m_wbs_dat_o_8[20] icon/m_wbs_dat_o_8[21] icon/m_wbs_dat_o_8[22]
+ icon/m_wbs_dat_o_8[23] icon/m_wbs_dat_o_8[24] icon/m_wbs_dat_o_8[25] icon/m_wbs_dat_o_8[26]
+ icon/m_wbs_dat_o_8[27] icon/m_wbs_dat_o_8[28] icon/m_wbs_dat_o_8[29] icon/m_wbs_dat_o_8[2]
+ icon/m_wbs_dat_o_8[30] icon/m_wbs_dat_o_8[31] icon/m_wbs_dat_o_8[3] icon/m_wbs_dat_o_8[4]
+ icon/m_wbs_dat_o_8[5] icon/m_wbs_dat_o_8[6] icon/m_wbs_dat_o_8[7] icon/m_wbs_dat_o_8[8]
+ icon/m_wbs_dat_o_8[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[8]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_7 wb_clk_i icon/m_wb_rst_i[7] icon/m_wbs_ack_o[7] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_7[0] icon/m_wbs_dat_o_7[10] icon/m_wbs_dat_o_7[11]
+ icon/m_wbs_dat_o_7[12] icon/m_wbs_dat_o_7[13] icon/m_wbs_dat_o_7[14] icon/m_wbs_dat_o_7[15]
+ icon/m_wbs_dat_o_7[16] icon/m_wbs_dat_o_7[17] icon/m_wbs_dat_o_7[18] icon/m_wbs_dat_o_7[19]
+ icon/m_wbs_dat_o_7[1] icon/m_wbs_dat_o_7[20] icon/m_wbs_dat_o_7[21] icon/m_wbs_dat_o_7[22]
+ icon/m_wbs_dat_o_7[23] icon/m_wbs_dat_o_7[24] icon/m_wbs_dat_o_7[25] icon/m_wbs_dat_o_7[26]
+ icon/m_wbs_dat_o_7[27] icon/m_wbs_dat_o_7[28] icon/m_wbs_dat_o_7[29] icon/m_wbs_dat_o_7[2]
+ icon/m_wbs_dat_o_7[30] icon/m_wbs_dat_o_7[31] icon/m_wbs_dat_o_7[3] icon/m_wbs_dat_o_7[4]
+ icon/m_wbs_dat_o_7[5] icon/m_wbs_dat_o_7[6] icon/m_wbs_dat_o_7[7] icon/m_wbs_dat_o_7[8]
+ icon/m_wbs_dat_o_7[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[7]
+ wbs_we_i vccd1 vssd1 ren_conv_top
Xren_conv_top_inst_9 wb_clk_i icon/m_wb_rst_i[9] icon/m_wbs_ack_o[9] wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] icon/m_wbs_dat_o_9[0] icon/m_wbs_dat_o_9[10] icon/m_wbs_dat_o_9[11]
+ icon/m_wbs_dat_o_9[12] icon/m_wbs_dat_o_9[13] icon/m_wbs_dat_o_9[14] icon/m_wbs_dat_o_9[15]
+ icon/m_wbs_dat_o_9[16] icon/m_wbs_dat_o_9[17] icon/m_wbs_dat_o_9[18] icon/m_wbs_dat_o_9[19]
+ icon/m_wbs_dat_o_9[1] icon/m_wbs_dat_o_9[20] icon/m_wbs_dat_o_9[21] icon/m_wbs_dat_o_9[22]
+ icon/m_wbs_dat_o_9[23] icon/m_wbs_dat_o_9[24] icon/m_wbs_dat_o_9[25] icon/m_wbs_dat_o_9[26]
+ icon/m_wbs_dat_o_9[27] icon/m_wbs_dat_o_9[28] icon/m_wbs_dat_o_9[29] icon/m_wbs_dat_o_9[2]
+ icon/m_wbs_dat_o_9[30] icon/m_wbs_dat_o_9[31] icon/m_wbs_dat_o_9[3] icon/m_wbs_dat_o_9[4]
+ icon/m_wbs_dat_o_9[5] icon/m_wbs_dat_o_9[6] icon/m_wbs_dat_o_9[7] icon/m_wbs_dat_o_9[8]
+ icon/m_wbs_dat_o_9[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] icon/m_wbs_stb_i[9]
+ wbs_we_i vccd1 vssd1 ren_conv_top
.ends

